VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_ef_ip__rc_osc_500k
  CLASS BLOCK ;
  FOREIGN sky130_ef_ip__rc_osc_500k ;
  ORIGIN 0.000 0.000 ;
  SIZE 61.210 BY 53.620 ;
  PIN avdd
    ANTENNADIFFAREA 148.754990 ;
    PORT
      LAYER met2 ;
        RECT -0.120 38.605 60.280 48.575 ;
    END
    PORT
      LAYER met2 ;
        RECT 60.720 38.605 61.220 48.575 ;
    END
  END avdd
  PIN avss
    ANTENNADIFFAREA 114.014595 ;
    PORT
      LAYER met2 ;
        RECT -0.120 5.250 1.595 15.220 ;
    END
    PORT
      LAYER met2 ;
        RECT 59.670 5.250 61.320 15.220 ;
    END
  END avss
  PIN dvss
    ANTENNADIFFAREA 6.628900 ;
    PORT
      LAYER met1 ;
        RECT 59.320 31.820 61.220 35.705 ;
    END
  END dvss
  PIN dvdd
    ANTENNADIFFAREA 4.280700 ;
    PORT
      LAYER met1 ;
        RECT 59.320 18.080 61.320 21.955 ;
    END
  END dvdd
  PIN ena
    ANTENNAGATEAREA 1.060500 ;
    ANTENNADIFFAREA 0.202500 ;
    PORT
      LAYER met2 ;
        RECT 60.210 23.930 61.210 24.930 ;
    END
  END ena
  PIN dout
    ANTENNADIFFAREA 0.556800 ;
    PORT
      LAYER met2 ;
        RECT 60.210 28.150 61.210 29.150 ;
    END
  END dout
  OBS
      LAYER nwell ;
        RECT -0.120 33.250 61.220 53.790 ;
        RECT -0.120 20.350 61.210 33.250 ;
        RECT -0.120 -0.190 61.320 20.350 ;
      LAYER li1 ;
        RECT 0.310 0.275 60.855 53.350 ;
      LAYER met1 ;
        RECT 0.310 35.985 60.770 51.100 ;
        RECT 0.310 31.540 59.040 35.985 ;
        RECT 0.310 22.235 60.770 31.540 ;
        RECT 0.310 17.800 59.040 22.235 ;
        RECT 0.310 2.490 60.770 17.800 ;
      LAYER met2 ;
        RECT 0.340 29.430 60.720 38.325 ;
        RECT 0.340 27.870 59.930 29.430 ;
        RECT 0.340 25.210 60.720 27.870 ;
        RECT 0.340 23.650 59.930 25.210 ;
        RECT 0.340 15.500 60.720 23.650 ;
        RECT 1.875 5.250 59.390 15.500 ;
      LAYER met3 ;
        RECT 11.160 13.590 37.435 28.385 ;
      LAYER met4 ;
        RECT 11.555 17.260 37.335 28.390 ;
  END
END sky130_ef_ip__rc_osc_500k
END LIBRARY

