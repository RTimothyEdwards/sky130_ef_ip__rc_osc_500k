* NGSPICE file created from sky130_ef_ip__rc_osc_500k.ext - technology: sky130A

.subckt sky130_ef_ip__rc_osc_500k dout ena dvss dvdd avdd avss
X0 a_1178_9768# a_1344_7168# avss.t90 sky130_fd_pr__res_xhigh_po_0p35 l=11
X1 a_10660_3118# a_10494_518# avss.t36 sky130_fd_pr__res_xhigh_po_0p35 l=11
X2 a_4352_3118# a_4186_518# avss.t148 sky130_fd_pr__res_xhigh_po_0p35 l=11
X3 a_6490_9768# a_6656_7168# avss.t85 sky130_fd_pr__res_xhigh_po_0p35 l=11
X4 a_3502_9768# a_3336_7168# avss.t0 sky130_fd_pr__res_xhigh_po_0p35 l=11
X5 a_5162_9768# a_4996_7168# avss.t159 sky130_fd_pr__res_xhigh_po_0p35 l=11
X6 a_8814_9768# a_8648_7168# avss.t119 sky130_fd_pr__res_xhigh_po_0p35 l=11
X7 a_2692_3118# a_2858_518# avss.t7 sky130_fd_pr__res_xhigh_po_0p35 l=11
X8 a_7718_4786# ena.t0 a_7560_4786# avss.t57 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X9 a_7154_9768# a_7320_7168# avss.t19 sky130_fd_pr__res_xhigh_po_0p35 l=11
X10 a_5348_3118# a_5182_518# avss.t87 sky130_fd_pr__res_xhigh_po_0p35 l=11
X11 a_11636_7168# a_11490_518# avss.t18 sky130_fd_pr__res_xhigh_po_0p35 l=11
X12 a_4166_9768# a_4000_7168# avss.t118 sky130_fd_pr__res_xhigh_po_0p35 l=11
X13 a_11138_9768# a_11304_7168# avss.t31 sky130_fd_pr__res_xhigh_po_0p35 l=11
X14 a_4194_4788.t1 a_3638_4788.t2 a_4036_4788# avss.t34 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X15 a_3688_3118# a_3854_518# avss.t101 sky130_fd_pr__res_xhigh_po_0p35 l=11
X16 a_2506_9768# a_2340_7168# avss.t43 sky130_fd_pr__res_xhigh_po_0p35 l=11
X17 a_9478_9768# a_9312_7168# avss.t29 sky130_fd_pr__res_xhigh_po_0p35 l=11
X18 a_7818_9768# a_7652_7168# avss.t62 sky130_fd_pr__res_xhigh_po_0p35 l=11
X19 a_6344_3118# a_6178_518# avss.t98 sky130_fd_pr__res_xhigh_po_0p35 l=11
X20 avdd.t16 a_2368_4788.t0 a_2368_4788.t1 avdd.t15 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X21 a_1032_3118# a_866_518# avss.t110 sky130_fd_pr__res_xhigh_po_0p35 l=11
X22 a_846_9768# a_1012_7168# avss.t54 sky130_fd_pr__res_xhigh_po_0p35 l=11
X23 a_6158_9768# a_6324_7168# avss.t111 sky130_fd_pr__res_xhigh_po_0p35 l=11
X24 a_4684_3118# a_4850_518# avss.t21 sky130_fd_pr__res_xhigh_po_0p35 l=11
X25 a_10806_9768# a_10972_7168# avss.t82 sky130_fd_pr__res_xhigh_po_0p35 l=11
X26 avss.t59 ena.t1 level_shifter_0.outb_h.t0 avss.t58 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X27 a_10142_9768# a_10308_7168# avss.t122 sky130_fd_pr__res_xhigh_po_0p35 l=11
X28 a_7340_3118# a_7174_518# avss.t24 sky130_fd_pr__res_xhigh_po_0p35 l=11
X29 avdd.t14 a_2368_4788.t4 a_4854_5653# avdd.t13 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X30 a_5826_9768# a_5992_7168# avss.t143 sky130_fd_pr__res_xhigh_po_0p35 l=11
X31 a_5162_9768# a_5328_7168# avss.t38 sky130_fd_pr__res_xhigh_po_0p35 l=11
X32 avdd.t12 a_2368_4788.t5 a_5470_5653# avdd.t11 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X33 a_2028_3118# a_1862_518# avss.t40 sky130_fd_pr__res_xhigh_po_0p35 l=11
X34 a_5680_3118# a_5846_518# avss.t23 sky130_fd_pr__res_xhigh_po_0p35 l=11
X35 a_9146_9768# a_8980_7168# avss.t1 sky130_fd_pr__res_xhigh_po_0p35 l=11
X36 a_8336_3118# a_8170_518# avss.t103 sky130_fd_pr__res_xhigh_po_0p35 l=11
X37 a_4830_9768# a_4996_7168# avss.t147 sky130_fd_pr__res_xhigh_po_0p35 l=11
X38 a_3024_3118# a_2858_518# avss.t146 sky130_fd_pr__res_xhigh_po_0p35 l=11
X39 a_6676_3118# a_6842_518# avss.t26 sky130_fd_pr__res_xhigh_po_0p35 l=11
X40 a_1364_3118# a_1530_518# avss.t131 sky130_fd_pr__res_xhigh_po_0p35 l=11
X41 a_10474_9768# a_10640_7168# avss.t56 sky130_fd_pr__res_xhigh_po_0p35 l=11
X42 a_1842_9768# a_1676_7168# avss.t30 sky130_fd_pr__res_xhigh_po_0p35 l=11
X43 a_9332_3118# a_9166_518# avss.t128 sky130_fd_pr__res_xhigh_po_0p35 l=11
X44 a_4020_3118# a_3854_518# avss.t125 sky130_fd_pr__res_xhigh_po_0p35 l=11
X45 avdd.t18 level_shifter_0.out_h.t2 a_2368_4788.t2 avdd.t15 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X46 a_3082_4788.t2 avss.t75 sky130_fd_pr__cap_mim_m3_1 l=6 w=3
X47 dvdd.t5 ena.t2 level_shifter_0.inb_l dvdd.t4 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X48 a_5494_9768# a_5660_7168# avss.t25 sky130_fd_pr__res_xhigh_po_0p35 l=11
X49 a_4750_4788.t1 a_4194_4788.t2 a_4854_5653# avdd.t13 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X50 a_10328_3118# a_10162_518# avss.t100 sky130_fd_pr__res_xhigh_po_0p35 l=11
X51 a_7672_3118# a_7838_518# avss.t112 sky130_fd_pr__res_xhigh_po_0p35 l=11
X52 a_1414_4786.t2 level_shifter_0.outb_h.t2 avss.t51 avss.t50 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X53 a_4750_4788.t2 avss.t86 sky130_fd_pr__cap_mim_m3_1 l=6 w=3
X54 a_700_3118# a_534_518# avss.t45 sky130_fd_pr__res_xhigh_po_0p35 l=11
X55 a_2360_3118# a_2526_518# avss.t107 sky130_fd_pr__res_xhigh_po_0p35 l=11
X56 a_1414_4786.t3 level_shifter_0.out_h.t3 a_514_7168# avss.t68 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X57 a_1032_3118# a_1198_518# avss.t124 sky130_fd_pr__res_xhigh_po_0p35 l=11
X58 a_3638_4788.t3 avss.t89 sky130_fd_pr__cap_mim_m3_1 l=6 w=3
X59 a_5306_4788.t1 a_4750_4788.t3 a_5470_5653# avdd.t11 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X60 a_11324_3118# a_11158_518# avss.t166 sky130_fd_pr__res_xhigh_po_0p35 l=11
X61 a_5016_3118# a_4850_518# avss.t66 sky130_fd_pr__res_xhigh_po_0p35 l=11
X62 a_4498_9768# a_4664_7168# avss.t11 sky130_fd_pr__res_xhigh_po_0p35 l=11
X63 a_8668_3118# a_8834_518# avss.t113 sky130_fd_pr__res_xhigh_po_0p35 l=11
X64 a_9810_9768# a_9976_7168# avss.t158 sky130_fd_pr__res_xhigh_po_0p35 l=11
X65 avdd.t10 a_2368_4788.t6 a_3622_5653# avdd.t9 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X66 a_3356_3118# a_3522_518# avss.t134 sky130_fd_pr__res_xhigh_po_0p35 l=11
X67 a_2028_3118# a_2194_518# avss.t102 sky130_fd_pr__res_xhigh_po_0p35 l=11
X68 a_6260_4788# a_1414_4786.t4 avss.t70 avss.t69 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X69 a_5306_4788.t2 avss.t149 sky130_fd_pr__cap_mim_m3_1 l=6 w=3
X70 a_3170_9768# a_3004_7168# avss.t164 sky130_fd_pr__res_xhigh_po_0p35 l=11
X71 a_6012_3118# a_5846_518# avss.t93 sky130_fd_pr__res_xhigh_po_0p35 l=11
X72 a_1510_9768# a_1344_7168# avss.t39 sky130_fd_pr__res_xhigh_po_0p35 l=11
X73 a_6822_9768# a_6656_7168# avss.t42 sky130_fd_pr__res_xhigh_po_0p35 l=11
X74 a_8482_9768# a_8316_7168# avss.t13 sky130_fd_pr__res_xhigh_po_0p35 l=11
X75 avdd.t8 a_2368_4788.t7 a_3006_5653# avdd.t7 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X76 a_9664_3118# a_9830_518# avss.t88 sky130_fd_pr__res_xhigh_po_0p35 l=11
X77 avdd.t6 a_2368_4788.t8 a_4238_5653# avdd.t5 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X78 dvss.t5 ena.t3 level_shifter_0.inb_l dvss.t4 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X79 a_10806_9768# a_10640_7168# avss.t14 sky130_fd_pr__res_xhigh_po_0p35 l=11
X80 a_9482_5327# level_shifter_0.out_h.t4 level_shifter_0.outb_h.t1 avdd.t21 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X81 a_3024_3118# a_3190_518# avss.t47 sky130_fd_pr__res_xhigh_po_0p35 l=11
X82 a_3502_9768# a_3668_7168# avss.t12 sky130_fd_pr__res_xhigh_po_0p35 l=11
X83 avdd.t4 a_2368_4788.t9 a_6702_5653# avdd.t3 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X84 a_4352_3118# a_4518_518# avss.t153 sky130_fd_pr__res_xhigh_po_0p35 l=11
X85 a_2174_9768# a_2008_7168# avss.t15 sky130_fd_pr__res_xhigh_po_0p35 l=11
X86 a_7486_9768# a_7320_7168# avss.t91 sky130_fd_pr__res_xhigh_po_0p35 l=11
X87 a_10660_3118# a_10826_518# avss.t77 sky130_fd_pr__res_xhigh_po_0p35 l=11
X88 a_5826_9768# a_5660_7168# avss.t126 sky130_fd_pr__res_xhigh_po_0p35 l=11
X89 dout.t0 a_7718_4786# dvdd.t1 dvdd.t0 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X90 a_7008_3118# a_6842_518# avss.t130 sky130_fd_pr__res_xhigh_po_0p35 l=11
X91 a_1696_3118# a_1530_518# avss.t117 sky130_fd_pr__res_xhigh_po_0p35 l=11
X92 avdd.t2 a_2368_4788.t10 a_6086_5653# avdd.t1 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X93 a_9332_3118# a_9498_518# avss.t133 sky130_fd_pr__res_xhigh_po_0p35 l=11
X94 a_11890_5939# a_7718_4786# dvss.t1 dvss.t0 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.15
D0 dvss.t3 ena.t4 sky130_fd_pr__diode_pw2nd_05v5 pj=1.8e+06 area=2.025e+11
X95 a_4166_9768# a_4332_7168# avss.t163 sky130_fd_pr__res_xhigh_po_0p35 l=11
X96 a_5348_3118# a_5514_518# avss.t129 sky130_fd_pr__res_xhigh_po_0p35 l=11
X97 a_4020_3118# a_4186_518# avss.t41 sky130_fd_pr__res_xhigh_po_0p35 l=11
X98 a_9478_9768# a_9644_7168# avss.t116 sky130_fd_pr__res_xhigh_po_0p35 l=11
X99 a_10328_3118# a_10494_518# avss.t115 sky130_fd_pr__res_xhigh_po_0p35 l=11
X100 a_514_9768# a_680_7168# avss.t156 sky130_fd_pr__res_xhigh_po_0p35 l=11
X101 level_shifter_0.out_h.t0 level_shifter_0.outb_h.t3 a_8714_4659# avdd.t17 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X102 a_1178_9768# a_1012_7168# avss.t22 sky130_fd_pr__res_xhigh_po_0p35 l=11
X103 a_8004_3118# a_7838_518# avss.t17 sky130_fd_pr__res_xhigh_po_0p35 l=11
X104 a_2692_3118# a_2526_518# avss.t27 sky130_fd_pr__res_xhigh_po_0p35 l=11
X105 a_5148_4788# a_1414_4786.t5 avss.t72 avss.t71 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X106 a_2982_4700.t0 a_5862_4788# a_6260_4788# avss.t69 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X107 a_8150_9768# a_7984_7168# avss.t76 sky130_fd_pr__res_xhigh_po_0p35 l=11
X108 level_shifter_0.out_h.t1 level_shifter_0.inb_l avss.t151 avss.t150 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X109 a_5704_4788# a_1414_4786.t6 avss.t73 avss.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X110 a_6344_3118# a_6510_518# avss.t20 sky130_fd_pr__res_xhigh_po_0p35 l=11
X111 a_3638_4788.t1 a_3082_4788.t3 a_3622_5653# avdd.t9 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X112 a_11324_3118# a_11490_518# avss.t120 sky130_fd_pr__res_xhigh_po_0p35 l=11
X113 a_5016_3118# a_5182_518# avss.t142 sky130_fd_pr__res_xhigh_po_0p35 l=11
X114 a_700_3118# a_866_518# avss.t127 sky130_fd_pr__res_xhigh_po_0p35 l=11
X115 a_9000_3118# a_8834_518# avss.t65 sky130_fd_pr__res_xhigh_po_0p35 l=11
X116 dvss.t7 level_shifter_0.inb_l dout.t2 dvss.t6 sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.15
X117 a_3480_4788# a_1414_4786.t7 avss.t74 avss.t52 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X118 a_3170_9768# a_3336_7168# avss.t28 sky130_fd_pr__res_xhigh_po_0p35 l=11
X119 a_8482_9768# a_8648_7168# avss.t104 sky130_fd_pr__res_xhigh_po_0p35 l=11
X120 a_3082_4788.t0 a_2982_4700.t2 a_3006_5653# avdd.t7 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X121 a_4194_4788.t0 a_3638_4788.t4 a_4238_5653# avdd.t5 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X122 dvdd.t3 ena.t5 a_7718_4786# dvdd.t2 sky130_fd_pr__pfet_01v8 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.15
X123 a_7154_9768# a_6988_7168# avss.t165 sky130_fd_pr__res_xhigh_po_0p35 l=11
X124 a_3688_3118# a_3522_518# avss.t63 sky130_fd_pr__res_xhigh_po_0p35 l=11
X125 a_11138_9768# a_10972_7168# avss.t99 sky130_fd_pr__res_xhigh_po_0p35 l=11
X126 a_2982_4700.t1 a_5862_4788# a_6702_5653# avdd.t3 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X127 a_7340_3118# a_7506_518# avss.t80 sky130_fd_pr__res_xhigh_po_0p35 l=11
X128 a_6012_3118# a_6178_518# avss.t135 sky130_fd_pr__res_xhigh_po_0p35 l=11
X129 a_3834_9768# a_4000_7168# avss.t136 sky130_fd_pr__res_xhigh_po_0p35 l=11
X130 a_9146_9768# a_9312_7168# avss.t81 sky130_fd_pr__res_xhigh_po_0p35 l=11
X131 a_9996_3118# a_9830_518# avss.t60 sky130_fd_pr__res_xhigh_po_0p35 l=11
X132 a_4684_3118# a_4518_518# avss.t132 sky130_fd_pr__res_xhigh_po_0p35 l=11
X133 a_5862_4788# a_5306_4788.t3 a_6086_5653# avdd.t1 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X134 a_10992_3118# a_10826_518# avss.t67 sky130_fd_pr__res_xhigh_po_0p35 l=11
X135 a_8336_3118# a_8502_518# avss.t61 sky130_fd_pr__res_xhigh_po_0p35 l=11
X136 a_6158_9768# a_5992_7168# avss.t94 sky130_fd_pr__res_xhigh_po_0p35 l=11
X137 a_5306_4788.t0 a_4750_4788.t4 a_5148_4788# avss.t71 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X138 a_7008_3118# a_7174_518# avss.t95 sky130_fd_pr__res_xhigh_po_0p35 l=11
X139 a_7718_4786# a_2982_4700.t3 dvdd.t6 avdd.t23 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X140 a_4592_4788# a_1414_4786.t8 avss.t137 avss.t5 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X141 a_5862_4788# a_5306_4788.t4 a_5704_4788# avss.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X142 a_846_9768# a_680_7168# avss.t32 sky130_fd_pr__res_xhigh_po_0p35 l=11
X143 a_8814_9768# a_8980_7168# avss.t161 sky130_fd_pr__res_xhigh_po_0p35 l=11
X144 a_5680_3118# a_5514_518# avss.t162 sky130_fd_pr__res_xhigh_po_0p35 l=11
X145 a_2838_9768# a_3004_7168# avss.t121 sky130_fd_pr__res_xhigh_po_0p35 l=11
X146 avdd.t22 level_shifter_0.out_h.t5 a_8714_4659# avdd.t17 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X147 a_8150_9768# a_8316_7168# avss.t96 sky130_fd_pr__res_xhigh_po_0p35 l=11
X148 a_3638_4788.t0 a_3082_4788.t4 a_3480_4788# avss.t52 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X149 a_2526_4188# a_1414_4786.t9 avss.t139 avss.t138 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X150 a_8004_3118# a_8170_518# avss.t33 sky130_fd_pr__res_xhigh_po_0p35 l=11
X151 a_2924_4788# a_1414_4786.t10 avss.t141 avss.t140 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X152 a_11470_9768# a_11304_7168# avss.t53 sky130_fd_pr__res_xhigh_po_0p35 l=11
X153 a_9482_5327# level_shifter_0.outb_h.t4 avdd.t20 avdd.t19 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X154 a_2506_9768# a_2672_7168# avss.t44 sky130_fd_pr__res_xhigh_po_0p35 l=11
X155 a_7818_9768# a_7984_7168# avss.t152 sky130_fd_pr__res_xhigh_po_0p35 l=11
X156 a_11890_5939# ena.t6 dout.t1 dvss.t2 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.15
X157 a_1842_9768# a_2008_7168# avss.t123 sky130_fd_pr__res_xhigh_po_0p35 l=11
X158 a_6676_3118# a_6510_518# avss.t10 sky130_fd_pr__res_xhigh_po_0p35 l=11
X159 a_6490_9768# a_6324_7168# avss.t3 sky130_fd_pr__res_xhigh_po_0p35 l=11
X160 a_1364_3118# a_1198_518# avss.t4 sky130_fd_pr__res_xhigh_po_0p35 l=11
X161 a_4830_9768# a_4664_7168# avss.t64 sky130_fd_pr__res_xhigh_po_0p35 l=11
X162 a_9000_3118# a_9166_518# avss.t108 sky130_fd_pr__res_xhigh_po_0p35 l=11
X163 a_10474_9768# a_10308_7168# avss.t109 sky130_fd_pr__res_xhigh_po_0p35 l=11
X164 a_9996_3118# a_10162_518# avss.t78 sky130_fd_pr__res_xhigh_po_0p35 l=11
X165 a_1510_9768# a_1676_7168# avss.t154 sky130_fd_pr__res_xhigh_po_0p35 l=11
X166 a_7672_3118# a_7506_518# avss.t155 sky130_fd_pr__res_xhigh_po_0p35 l=11
X167 a_514_9768# a_514_7168# avss.t97 sky130_fd_pr__res_xhigh_po_0p35 l=11
X168 a_6822_9768# a_6988_7168# avss.t9 sky130_fd_pr__res_xhigh_po_0p35 l=11
X169 a_4750_4788.t0 a_4194_4788.t3 a_4592_4788# avss.t5 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X170 a_2360_3118# a_2194_518# avss.t55 sky130_fd_pr__res_xhigh_po_0p35 l=11
X171 a_4194_4788.t4 avss.t6 sky130_fd_pr__cap_mim_m3_1 l=6 w=3
X172 a_5494_9768# a_5328_7168# avss.t114 sky130_fd_pr__res_xhigh_po_0p35 l=11
X173 a_2526_4188# level_shifter_0.out_h.t6 a_2368_4788.t3 avss.t138 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X174 a_3834_9768# a_3668_7168# avss.t49 sky130_fd_pr__res_xhigh_po_0p35 l=11
X175 a_3082_4788.t1 a_2982_4700.t4 a_2924_4788# avss.t140 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X176 avdd a_534_518# avss.t2 sky130_fd_pr__res_xhigh_po_0p35 l=11
X177 a_1414_4786.t1 a_1414_4786.t0 avss.t92 avss.t68 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X178 a_7560_4786# a_2982_4700.t5 avss.t160 avss.t57 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X179 a_2174_9768# a_2340_7168# avss.t46 sky130_fd_pr__res_xhigh_po_0p35 l=11
X180 a_7486_9768# a_7652_7168# avss.t83 sky130_fd_pr__res_xhigh_po_0p35 l=11
X181 a_10992_3118# a_11158_518# avss.t84 sky130_fd_pr__res_xhigh_po_0p35 l=11
X182 a_8668_3118# a_8502_518# avss.t79 sky130_fd_pr__res_xhigh_po_0p35 l=11
X183 a_3356_3118# a_3190_518# avss.t37 sky130_fd_pr__res_xhigh_po_0p35 l=11
X184 a_4036_4788# a_1414_4786.t11 avss.t35 avss.t34 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X185 a_11470_9768# a_11636_7168# avss.t105 sky130_fd_pr__res_xhigh_po_0p35 l=11
X186 a_2838_9768# a_2672_7168# avss.t106 sky130_fd_pr__res_xhigh_po_0p35 l=11
X187 a_4498_9768# a_4332_7168# avss.t48 sky130_fd_pr__res_xhigh_po_0p35 l=11
X188 a_9810_9768# a_9644_7168# avss.t144 sky130_fd_pr__res_xhigh_po_0p35 l=11
X189 a_1696_3118# a_1862_518# avss.t145 sky130_fd_pr__res_xhigh_po_0p35 l=11
X190 a_9664_3118# a_9498_518# avss.t8 sky130_fd_pr__res_xhigh_po_0p35 l=11
X191 a_10142_9768# a_9976_7168# avss.t157 sky130_fd_pr__res_xhigh_po_0p35 l=11
R0 avss.n269 avss.n3 42418.7
R1 avss.n348 avss.n3 42418.7
R2 avss.n348 avss.n4 42418.7
R3 avss.n269 avss.n4 42418.7
R4 avss.n36 avss.n28 42418.7
R5 avss.n322 avss.n28 42418.7
R6 avss.n322 avss.n29 42418.7
R7 avss.n36 avss.n29 42418.7
R8 avss.n300 avss.n299 4540.48
R9 avss.n324 avss.n323 3194
R10 avss.n301 avss.n39 1379.81
R11 avss.n301 avss.n40 1379.81
R12 avss.n314 avss.n40 1379.81
R13 avss.n314 avss.n39 1379.81
R14 avss.n346 avss.n5 1379.81
R15 avss.n346 avss.n6 1379.81
R16 avss.n326 avss.n6 1379.81
R17 avss.n326 avss.n5 1379.81
R18 avss.n331 avss.n22 1379.81
R19 avss.n332 avss.n22 1379.81
R20 avss.n332 avss.n21 1379.81
R21 avss.n331 avss.n21 1379.81
R22 avss.n215 avss.n214 1379.81
R23 avss.n220 avss.n215 1379.81
R24 avss.n221 avss.n220 1379.81
R25 avss.n221 avss.n214 1379.81
R26 avss.n235 avss.n105 1379.81
R27 avss.n234 avss.n105 1379.81
R28 avss.n234 avss.n104 1379.81
R29 avss.n235 avss.n104 1379.81
R30 avss.n240 avss.n98 1379.81
R31 avss.n241 avss.n98 1379.81
R32 avss.n241 avss.n97 1379.81
R33 avss.n240 avss.n97 1379.81
R34 avss.n189 avss.n182 1379.81
R35 avss.n182 avss.n123 1379.81
R36 avss.n178 avss.n123 1379.81
R37 avss.n189 avss.n178 1379.81
R38 avss.n253 avss.n81 1379.81
R39 avss.n252 avss.n81 1379.81
R40 avss.n252 avss.n80 1379.81
R41 avss.n253 avss.n80 1379.81
R42 avss.n258 avss.n74 1379.81
R43 avss.n259 avss.n74 1379.81
R44 avss.n259 avss.n73 1379.81
R45 avss.n258 avss.n73 1379.81
R46 avss.n162 avss.n140 1379.81
R47 avss.n140 avss.n135 1379.81
R48 avss.n136 avss.n135 1379.81
R49 avss.n162 avss.n136 1379.81
R50 avss.n156 avss.n57 1379.81
R51 avss.n156 avss.n58 1379.81
R52 avss.n288 avss.n58 1379.81
R53 avss.n288 avss.n57 1379.81
R54 avss.n290 avss.n49 1379.81
R55 avss.n290 avss.n50 1379.81
R56 avss.n297 avss.n50 1379.81
R57 avss.n297 avss.n49 1379.81
R58 avss.n202 avss.n18 1379.81
R59 avss.n202 avss.n23 1379.81
R60 avss.n217 avss.n23 1379.81
R61 avss.n217 avss.n18 1379.81
R62 avss.n216 avss.n200 1379.81
R63 avss.n216 avss.n208 1379.81
R64 avss.n223 avss.n208 1379.81
R65 avss.n223 avss.n200 1379.81
R66 avss.n209 avss.n106 1379.81
R67 avss.n209 avss.n107 1379.81
R68 avss.n114 avss.n107 1379.81
R69 avss.n114 avss.n106 1379.81
R70 avss.n117 avss.n95 1379.81
R71 avss.n117 avss.n99 1379.81
R72 avss.n179 avss.n99 1379.81
R73 avss.n179 avss.n95 1379.81
R74 avss.n122 avss.n121 1379.81
R75 avss.n190 avss.n121 1379.81
R76 avss.n190 avss.n120 1379.81
R77 avss.n122 avss.n120 1379.81
R78 avss.n175 avss.n82 1379.81
R79 avss.n175 avss.n83 1379.81
R80 avss.n126 avss.n83 1379.81
R81 avss.n126 avss.n82 1379.81
R82 avss.n129 avss.n71 1379.81
R83 avss.n129 avss.n75 1379.81
R84 avss.n137 avss.n75 1379.81
R85 avss.n137 avss.n71 1379.81
R86 avss.n134 avss.n133 1379.81
R87 avss.n163 avss.n133 1379.81
R88 avss.n163 avss.n132 1379.81
R89 avss.n134 avss.n132 1379.81
R90 avss.n152 avss.n62 1379.81
R91 avss.n152 avss.n144 1379.81
R92 avss.n144 avss.n56 1379.81
R93 avss.n62 avss.n56 1379.81
R94 avss.n292 avss.n54 1379.81
R95 avss.n55 avss.n54 1379.81
R96 avss.n55 avss.n48 1379.81
R97 avss.n292 avss.n48 1379.81
R98 avss.n308 avss.n45 1379.81
R99 avss.n310 avss.n44 1379.81
R100 avss.n310 avss.n45 1379.81
R101 avss.t58 avss.n35 934.398
R102 avss.n300 avss.t150 934.398
R103 avss.n321 avss.n30 812.683
R104 avss.n270 avss.n2 804.212
R105 avss.n349 avss.n2 800.46
R106 avss.n31 avss.n30 789.457
R107 avss.n315 avss.n38 697.509
R108 avss.n321 avss.n320 691.125
R109 avss.n271 avss.n268 665.563
R110 avss.n309 avss.n44 562.854
R111 avss.n316 avss.n35 552.742
R112 avss.n319 avss.n31 460.964
R113 avss.n350 avss.n1 360.981
R114 avss.n320 avss.n319 326.962
R115 avss.n267 avss.n1 307.827
R116 avss.n316 avss.n315 236.889
R117 avss.t150 avss.n38 236.889
R118 avss.n64 avss.t160 235.553
R119 avss.n343 avss.t51 234.381
R120 avss.n283 avss.t70 234.012
R121 avss.n264 avss.t73 234.012
R122 avss.n87 avss.t72 234.012
R123 avss.n249 avss.t137 234.012
R124 avss.n246 avss.t35 234.012
R125 avss.n227 avss.t74 234.012
R126 avss.n231 avss.t141 234.012
R127 avss.n337 avss.t139 234.012
R128 avss.n19 avss.t92 233.994
R129 avss.n46 avss.t59 233.939
R130 avss.n33 avss.t151 233.929
R131 avss.t18 avss.t120 213.194
R132 avss.t120 avss.t166 213.194
R133 avss.t166 avss.t84 213.194
R134 avss.t84 avss.t67 213.194
R135 avss.t67 avss.t77 213.194
R136 avss.t77 avss.t36 213.194
R137 avss.t36 avss.t115 213.194
R138 avss.t115 avss.t100 213.194
R139 avss.t100 avss.t78 213.194
R140 avss.t78 avss.t60 213.194
R141 avss.t60 avss.t88 213.194
R142 avss.t53 avss.t105 212.946
R143 avss.t31 avss.t53 212.946
R144 avss.t99 avss.t31 212.946
R145 avss.t82 avss.t99 212.946
R146 avss.t14 avss.t82 212.946
R147 avss.t56 avss.t14 212.946
R148 avss.t109 avss.t56 212.946
R149 avss.t122 avss.t109 212.946
R150 avss.t157 avss.t122 212.946
R151 avss.t158 avss.t157 212.946
R152 avss.t144 avss.t158 212.946
R153 avss.t116 avss.t144 204.929
R154 avss.t88 avss.t8 204.137
R155 avss.n269 avss.t18 202.793
R156 avss.t105 avss.n36 202.572
R157 avss.t29 avss.t116 197.994
R158 avss.t81 avss.t29 197.994
R159 avss.t1 avss.t81 197.994
R160 avss.t161 avss.t1 197.994
R161 avss.t119 avss.t104 197.994
R162 avss.t104 avss.t13 197.994
R163 avss.t13 avss.t96 197.994
R164 avss.t96 avss.t76 197.994
R165 avss.t76 avss.t152 197.994
R166 avss.t152 avss.t62 197.994
R167 avss.t62 avss.t83 197.994
R168 avss.t83 avss.t91 197.994
R169 avss.t91 avss.t19 197.994
R170 avss.t19 avss.t165 197.994
R171 avss.t165 avss.t9 197.964
R172 avss.t9 avss.t42 197.94
R173 avss.t42 avss.t85 197.94
R174 avss.t85 avss.t3 197.94
R175 avss.t3 avss.t111 197.94
R176 avss.t111 avss.t94 197.94
R177 avss.t143 avss.t126 197.94
R178 avss.t126 avss.t25 197.94
R179 avss.t25 avss.t114 197.94
R180 avss.t114 avss.t38 197.94
R181 avss.t38 avss.t159 197.94
R182 avss.t159 avss.t147 197.94
R183 avss.t147 avss.t64 197.94
R184 avss.t64 avss.t11 197.94
R185 avss.t11 avss.t48 197.94
R186 avss.t48 avss.t163 197.94
R187 avss.t163 avss.t118 197.94
R188 avss.t118 avss.t136 197.94
R189 avss.t136 avss.t49 197.94
R190 avss.t49 avss.t12 197.94
R191 avss.t12 avss.t0 197.94
R192 avss.t0 avss.t28 197.94
R193 avss.t28 avss.t164 197.94
R194 avss.t164 avss.t121 197.94
R195 avss.t121 avss.t106 197.94
R196 avss.t106 avss.t44 197.94
R197 avss.t44 avss.t43 197.94
R198 avss.t43 avss.t46 197.94
R199 avss.t46 avss.t15 197.94
R200 avss.t15 avss.t123 197.94
R201 avss.t123 avss.t30 197.94
R202 avss.t30 avss.t154 197.94
R203 avss.t154 avss.t39 197.94
R204 avss.t39 avss.t90 197.94
R205 avss.t22 avss.t54 197.94
R206 avss.t54 avss.t32 197.94
R207 avss.t32 avss.t156 197.94
R208 avss.t156 avss.t97 197.94
R209 avss.t8 avss.t133 191.405
R210 avss.t133 avss.t128 191.405
R211 avss.t128 avss.t108 191.405
R212 avss.t108 avss.t65 191.405
R213 avss.t65 avss.t113 191.405
R214 avss.t113 avss.t79 191.405
R215 avss.t79 avss.t61 191.405
R216 avss.t97 avss.n322 189.195
R217 avss.n38 avss.t161 163.405
R218 avss.n323 avss.t90 146.667
R219 avss.n293 avss.n292 146.25
R220 avss.n292 avss.t57 146.25
R221 avss.n146 avss.n55 146.25
R222 avss.t57 avss.n55 146.25
R223 avss.n285 avss.n62 146.25
R224 avss.t69 avss.n62 146.25
R225 avss.n149 avss.n144 146.25
R226 avss.n144 avss.t69 146.25
R227 avss.n134 avss.n66 146.25
R228 avss.t16 avss.n134 146.25
R229 avss.n164 avss.n163 146.25
R230 avss.n163 avss.t16 146.25
R231 avss.n260 avss.n71 146.25
R232 avss.t71 avss.n71 146.25
R233 avss.n167 avss.n75 146.25
R234 avss.t71 avss.n75 146.25
R235 avss.n251 avss.n82 146.25
R236 avss.t5 avss.n82 146.25
R237 avss.n170 avss.n83 146.25
R238 avss.t5 avss.n83 146.25
R239 avss.n122 avss.n90 146.25
R240 avss.t34 avss.n122 146.25
R241 avss.n191 avss.n190 146.25
R242 avss.n190 avss.t34 146.25
R243 avss.n242 avss.n95 146.25
R244 avss.t52 avss.n95 146.25
R245 avss.n194 avss.n99 146.25
R246 avss.t52 avss.n99 146.25
R247 avss.n233 avss.n106 146.25
R248 avss.t140 avss.n106 146.25
R249 avss.n197 avss.n107 146.25
R250 avss.t140 avss.n107 146.25
R251 avss.n200 avss.n13 146.25
R252 avss.t138 avss.n200 146.25
R253 avss.n208 avss.n207 146.25
R254 avss.t138 avss.n208 146.25
R255 avss.n333 avss.n18 146.25
R256 avss.t68 avss.n18 146.25
R257 avss.n204 avss.n23 146.25
R258 avss.t68 avss.n23 146.25
R259 avss.n295 avss.n49 146.25
R260 avss.t57 avss.n49 146.25
R261 avss.n293 avss.n50 146.25
R262 avss.t57 avss.n50 146.25
R263 avss.n61 avss.n57 146.25
R264 avss.t69 avss.n57 146.25
R265 avss.n285 avss.n58 146.25
R266 avss.t69 avss.n58 146.25
R267 avss.n162 avss.n161 146.25
R268 avss.t16 avss.n162 146.25
R269 avss.n135 avss.n66 146.25
R270 avss.t16 avss.n135 146.25
R271 avss.n258 avss.n257 146.25
R272 avss.t71 avss.n258 146.25
R273 avss.n260 avss.n259 146.25
R274 avss.n259 avss.t71 146.25
R275 avss.n254 avss.n253 146.25
R276 avss.n253 avss.t5 146.25
R277 avss.n252 avss.n251 146.25
R278 avss.t5 avss.n252 146.25
R279 avss.n189 avss.n188 146.25
R280 avss.t34 avss.n189 146.25
R281 avss.n123 avss.n90 146.25
R282 avss.t34 avss.n123 146.25
R283 avss.n240 avss.n239 146.25
R284 avss.t52 avss.n240 146.25
R285 avss.n242 avss.n241 146.25
R286 avss.n241 avss.t52 146.25
R287 avss.n236 avss.n235 146.25
R288 avss.n235 avss.t140 146.25
R289 avss.n234 avss.n233 146.25
R290 avss.t140 avss.n234 146.25
R291 avss.n214 avss.n213 146.25
R292 avss.t138 avss.n214 146.25
R293 avss.n220 avss.n13 146.25
R294 avss.n220 avss.t138 146.25
R295 avss.n331 avss.n330 146.25
R296 avss.t68 avss.n331 146.25
R297 avss.n333 avss.n332 146.25
R298 avss.n332 avss.t68 146.25
R299 avss.n7 avss.n5 146.25
R300 avss.t50 avss.n5 146.25
R301 avss.n8 avss.n6 146.25
R302 avss.t50 avss.n6 146.25
R303 avss.n304 avss.n39 146.25
R304 avss.t150 avss.n39 146.25
R305 avss.n42 avss.n40 146.25
R306 avss.t150 avss.n40 146.25
R307 avss.n311 avss.n310 146.25
R308 avss.n310 avss.t58 146.25
R309 avss.n308 avss.n307 146.25
R310 avss.t33 avss.t17 145.094
R311 avss.t155 avss.t112 145.094
R312 avss.t24 avss.t95 145.094
R313 avss.t95 avss.t130 145.094
R314 avss.t130 avss.t26 145.094
R315 avss.t26 avss.t10 145.094
R316 avss.t98 avss.t20 145.094
R317 avss.t66 avss.t142 145.094
R318 avss.t21 avss.t132 145.094
R319 avss.t37 avss.t134 145.094
R320 avss.t47 avss.t146 145.094
R321 avss.t117 avss.t145 145.094
R322 avss.t131 avss.t4 145.094
R323 avss.t127 avss.t110 145.094
R324 avss.t45 avss.t127 145.094
R325 avss.t2 avss.t45 145.094
R326 avss.n348 avss.t2 142.078
R327 avss.t17 avss.n298 138.101
R328 avss.t61 avss.t103 136.425
R329 avss.t69 avss.t135 135.48
R330 avss.t5 avss.t153 128.487
R331 avss.n153 avss.t23 125.865
R332 avss.t68 avss.t40 124.99
R333 avss.t140 avss.t7 121.495
R334 avss.n177 avss.t41 118.873
R335 avss.t52 avss.t63 117.999
R336 avss.n145 avss.n48 117.207
R337 avss.n298 avss.n48 117.001
R338 avss.n54 avss.n52 117.001
R339 avss.n291 avss.n54 117.001
R340 avss.n59 avss.n56 117.001
R341 avss.n289 avss.n56 117.001
R342 avss.n152 avss.n151 117.001
R343 avss.n155 avss.n152 117.001
R344 avss.n141 avss.n132 117.001
R345 avss.n153 avss.n132 117.001
R346 avss.n133 avss.n68 117.001
R347 avss.n139 avss.n133 117.001
R348 avss.n137 avss.n70 117.001
R349 avss.n138 avss.n137 117.001
R350 avss.n130 avss.n129 117.001
R351 avss.n129 avss.n128 117.001
R352 avss.n126 avss.n124 117.001
R353 avss.n127 avss.n126 117.001
R354 avss.n175 avss.n174 117.001
R355 avss.n176 avss.n175 117.001
R356 avss.n183 avss.n120 117.001
R357 avss.n177 avss.n120 117.001
R358 avss.n121 avss.n92 117.001
R359 avss.n181 avss.n121 117.001
R360 avss.n179 avss.n94 117.001
R361 avss.n180 avss.n179 117.001
R362 avss.n118 avss.n117 117.001
R363 avss.n117 avss.n116 117.001
R364 avss.n114 avss.n112 117.001
R365 avss.n115 avss.n114 117.001
R366 avss.n209 avss.n110 117.001
R367 avss.n210 avss.n209 117.001
R368 avss.n224 avss.n223 117.001
R369 avss.n223 avss.n222 117.001
R370 avss.n216 avss.n15 117.001
R371 avss.n219 avss.n216 117.001
R372 avss.n217 avss.n17 117.001
R373 avss.n218 avss.n217 117.001
R374 avss.n203 avss.n202 117.001
R375 avss.n202 avss.n27 117.001
R376 avss.n297 avss.n296 117.001
R377 avss.n298 avss.n297 117.001
R378 avss.n290 avss.n53 117.001
R379 avss.n291 avss.n290 117.001
R380 avss.n288 avss.n287 117.001
R381 avss.n289 avss.n288 117.001
R382 avss.n157 avss.n156 117.001
R383 avss.n156 avss.n155 117.001
R384 avss.n143 avss.n136 117.001
R385 avss.n153 avss.n136 117.001
R386 avss.n140 avss.n67 117.001
R387 avss.n140 avss.n139 117.001
R388 avss.n73 avss.n69 117.001
R389 avss.n138 avss.n73 117.001
R390 avss.n77 avss.n74 117.001
R391 avss.n128 avss.n74 117.001
R392 avss.n80 avss.n78 117.001
R393 avss.n127 avss.n80 117.001
R394 avss.n85 avss.n81 117.001
R395 avss.n176 avss.n81 117.001
R396 avss.n185 avss.n178 117.001
R397 avss.n178 avss.n177 117.001
R398 avss.n182 avss.n91 117.001
R399 avss.n182 avss.n181 117.001
R400 avss.n97 avss.n93 117.001
R401 avss.n180 avss.n97 117.001
R402 avss.n101 avss.n98 117.001
R403 avss.n116 avss.n98 117.001
R404 avss.n104 avss.n102 117.001
R405 avss.n115 avss.n104 117.001
R406 avss.n109 avss.n105 117.001
R407 avss.n210 avss.n105 117.001
R408 avss.n221 avss.n111 117.001
R409 avss.n222 avss.n221 117.001
R410 avss.n215 avss.n14 117.001
R411 avss.n219 avss.n215 117.001
R412 avss.n21 avss.n16 117.001
R413 avss.n218 avss.n21 117.001
R414 avss.n25 avss.n22 117.001
R415 avss.n27 avss.n22 117.001
R416 avss.n327 avss.n326 117.001
R417 avss.n326 avss.n325 117.001
R418 avss.n346 avss.n345 117.001
R419 avss.n347 avss.n346 117.001
R420 avss.n302 avss.n301 117.001
R421 avss.n301 avss.n300 117.001
R422 avss.n45 avss.n41 117.001
R423 avss.n45 avss.n35 117.001
R424 avss.n314 avss.n313 117.001
R425 avss.n315 avss.n314 117.001
R426 avss.n44 avss.n43 117.001
R427 avss.t55 avss.n219 115.376
R428 avss.t10 avss.n289 113.627
R429 avss.n128 avss.n127 113.627
R430 avss.n116 avss.n115 113.627
R431 avss.n325 avss.n27 113.627
R432 avss.n222 avss.t107 111.879
R433 avss.t57 avss.t80 111.005
R434 avss.t71 avss.t87 111.005
R435 avss.n181 avss.t125 108.383
R436 avss.n299 avss.t103 104.888
R437 avss.n139 avss.t162 101.391
R438 avss.t94 avss.n37 98.9707
R439 avss.n37 avss.t143 98.9707
R440 avss.n204 avss.n203 98.8418
R441 avss.t50 avss.n324 94.3986
R442 avss.t148 avss.n176 87.4061
R443 avss.t16 avss.t162 84.784
R444 avss.t102 avss.n218 83.9099
R445 avss.n294 avss.n52 82.4476
R446 avss.n287 avss.n59 82.0711
R447 avss.n328 avss.n327 82.0711
R448 avss.n327 avss.n26 82.0711
R449 avss.n151 avss.n63 82.0711
R450 avss.n225 avss.n111 82.0711
R451 avss.n225 avss.n224 82.0711
R452 avss.n335 avss.n14 82.0711
R453 avss.n335 avss.n15 82.0711
R454 avss.n108 avss.n102 82.0711
R455 avss.n112 avss.n108 82.0711
R456 avss.n226 avss.n109 82.0711
R457 avss.n226 avss.n110 82.0711
R458 avss.n243 avss.n93 82.0711
R459 avss.n243 avss.n94 82.0711
R460 avss.n113 avss.n101 82.0711
R461 avss.n118 avss.n113 82.0711
R462 avss.n185 avss.n184 82.0711
R463 avss.n184 avss.n183 82.0711
R464 avss.n244 avss.n91 82.0711
R465 avss.n244 avss.n92 82.0711
R466 avss.n84 avss.n78 82.0711
R467 avss.n124 avss.n84 82.0711
R468 avss.n86 avss.n85 82.0711
R469 avss.n174 avss.n86 82.0711
R470 avss.n261 avss.n69 82.0711
R471 avss.n261 avss.n70 82.0711
R472 avss.n125 avss.n77 82.0711
R473 avss.n130 avss.n125 82.0711
R474 avss.n143 avss.n142 82.0711
R475 avss.n142 avss.n141 82.0711
R476 avss.n262 avss.n67 82.0711
R477 avss.n262 avss.n68 82.0711
R478 avss.n157 avss.n63 82.0711
R479 avss.n329 avss.n25 82.0711
R480 avss.n201 avss.n25 82.0711
R481 avss.n24 avss.n16 82.0711
R482 avss.n334 avss.n16 82.0711
R483 avss.n334 avss.n17 82.0711
R484 avss.n203 avss.n201 82.0711
R485 avss.n148 avss.n59 81.6946
R486 avss.n151 avss.n150 81.6946
R487 avss.n211 avss.n111 81.6946
R488 avss.n224 avss.n199 81.6946
R489 avss.n212 avss.n14 81.6946
R490 avss.n206 avss.n15 81.6946
R491 avss.n237 avss.n102 81.6946
R492 avss.n196 avss.n112 81.6946
R493 avss.n109 avss.n103 81.6946
R494 avss.n198 avss.n110 81.6946
R495 avss.n100 avss.n93 81.6946
R496 avss.n193 avss.n94 81.6946
R497 avss.n238 avss.n101 81.6946
R498 avss.n195 avss.n118 81.6946
R499 avss.n186 avss.n185 81.6946
R500 avss.n183 avss.n119 81.6946
R501 avss.n187 avss.n91 81.6946
R502 avss.n192 avss.n92 81.6946
R503 avss.n255 avss.n78 81.6946
R504 avss.n169 avss.n124 81.6946
R505 avss.n85 avss.n79 81.6946
R506 avss.n174 avss.n173 81.6946
R507 avss.n76 avss.n69 81.6946
R508 avss.n166 avss.n70 81.6946
R509 avss.n256 avss.n77 81.6946
R510 avss.n168 avss.n130 81.6946
R511 avss.n159 avss.n143 81.6946
R512 avss.n141 avss.n131 81.6946
R513 avss.n160 avss.n67 81.6946
R514 avss.n165 avss.n68 81.6946
R515 avss.n158 avss.n157 81.6946
R516 avss.n205 avss.n17 81.6946
R517 avss.n147 avss.n52 80.9417
R518 avss.t27 avss.n210 80.4137
R519 avss.n309 avss.n308 78.2942
R520 avss.t34 avss.t125 77.7915
R521 avss.t101 avss.n180 76.9175
R522 avss.n317 avss.n316 75.7785
R523 avss.t80 avss.n291 75.1694
R524 avss.n138 avss.t87 75.1694
R525 avss.t138 avss.t107 74.2953
R526 avss.t110 avss.n347 73.4212
R527 avss.n154 avss.t93 72.5472
R528 avss.n347 avss.t124 71.6731
R529 avss.t138 avss.t55 70.7991
R530 avss.n148 avss.n147 70.3602
R531 avss.n291 avss.t24 69.925
R532 avss.t129 avss.n138 69.925
R533 avss.n180 avss.t63 68.1769
R534 avss.t34 avss.t41 67.3028
R535 avss.n210 avss.t7 64.6807
R536 avss.n218 avss.t40 61.1844
R537 avss.t16 avss.t23 60.3104
R538 avss.t58 avss.n309 59.6593
R539 avss.n176 avss.t153 57.6882
R540 avss.n323 avss.t22 51.2742
R541 avss.n155 avss.t135 50.6958
R542 avss.n311 avss.n43 50.3092
R543 avss.n302 avss.n42 50.106
R544 avss.n139 avss.t129 43.7033
R545 avss.n296 avss.n295 43.1857
R546 avss.n345 avss.n7 41.347
R547 avss.n303 avss.n302 40.4775
R548 avss.n299 avss.t33 40.2071
R549 avss.n146 avss.n145 39.9597
R550 avss.n47 avss.n43 39.8117
R551 avss.n181 avss.t101 36.7109
R552 avss.n38 avss.t119 34.5898
R553 avss.t57 avss.t155 34.0887
R554 avss.t71 avss.t142 34.0887
R555 avss.n222 avss.t27 33.2146
R556 avss.n289 avss.t20 31.4665
R557 avss.t4 avss.t50 30.5925
R558 avss.n219 avss.t102 29.7184
R559 avss.n345 avss.n344 27.9126
R560 avss.t52 avss.t134 27.0962
R561 avss.n177 avss.t148 26.2222
R562 avss.n145 avss.n51 25.3701
R563 avss.n296 avss.n51 25.361
R564 avss.n127 avss.t21 24.4741
R565 avss.n312 avss.n311 23.6684
R566 avss.t140 avss.t146 23.6
R567 avss.n312 avss.n42 23.4269
R568 avss.n155 avss.n154 21.8519
R569 avss.n27 avss.t117 20.9779
R570 avss.t68 avss.t145 20.1038
R571 avss.n324 avss.t124 20.1038
R572 avss.t93 avss.n153 19.2297
R573 avss.n293 avss.n51 17.4857
R574 avss.n115 avss.t47 17.4816
R575 avss.n158 avss.n61 17.1477
R576 avss.n161 avss.n159 17.1477
R577 avss.n161 avss.n160 17.1477
R578 avss.n257 avss.n76 17.1477
R579 avss.n257 avss.n256 17.1477
R580 avss.n255 avss.n254 17.1477
R581 avss.n254 avss.n79 17.1477
R582 avss.n188 avss.n186 17.1477
R583 avss.n188 avss.n187 17.1477
R584 avss.n239 avss.n100 17.1477
R585 avss.n239 avss.n238 17.1477
R586 avss.n237 avss.n236 17.1477
R587 avss.n236 avss.n103 17.1477
R588 avss.n213 avss.n211 17.1477
R589 avss.n213 avss.n212 17.1477
R590 avss.n147 avss.n146 17.1477
R591 avss.n149 avss.n148 17.1477
R592 avss.n150 avss.n149 17.1477
R593 avss.n164 avss.n131 17.1477
R594 avss.n165 avss.n164 17.1477
R595 avss.n167 avss.n166 17.1477
R596 avss.n168 avss.n167 17.1477
R597 avss.n170 avss.n169 17.1477
R598 avss.n191 avss.n119 17.1477
R599 avss.n192 avss.n191 17.1477
R600 avss.n194 avss.n193 17.1477
R601 avss.n195 avss.n194 17.1477
R602 avss.n197 avss.n196 17.1477
R603 avss.n198 avss.n197 17.1477
R604 avss.n207 avss.n199 17.1477
R605 avss.n207 avss.n206 17.1477
R606 avss.n205 avss.n204 17.1477
R607 avss.n328 avss.n7 17.0405
R608 avss.n330 avss.n24 17.0405
R609 avss.n330 avss.n329 17.0405
R610 avss.n26 avss.n8 16.8301
R611 avss.n334 avss.n333 16.8301
R612 avss.n225 avss.n13 16.6249
R613 avss.n233 avss.n108 16.6249
R614 avss.n243 avss.n242 16.6249
R615 avss.n184 avss.n90 16.6249
R616 avss.n251 avss.n84 16.6249
R617 avss.n261 avss.n260 16.6249
R618 avss.n142 avss.n66 16.6249
R619 avss.t5 avss.t132 16.6076
R620 avss.n286 avss.n61 15.7791
R621 avss.n313 avss.n312 15.7042
R622 avss.n295 avss.n294 15.6805
R623 avss.n286 avss.n285 15.2981
R624 avss.n294 avss.n293 15.2981
R625 avss.n307 avss.n306 15.1138
R626 avss.n306 avss.n304 14.9595
R627 avss.n172 avss.n170 14.4911
R628 avss.n116 avss.t37 13.9854
R629 avss.n305 avss.n41 13.6894
R630 avss.n270 avss.n269 12.7179
R631 avss.n36 avss.n31 12.7179
R632 avss.n322 avss.n321 12.7179
R633 avss.n349 avss.n348 12.7179
R634 avss.n344 avss.n8 12.7033
R635 avss.n325 avss.t131 10.4892
R636 avss.n159 avss.n158 10.4659
R637 avss.n160 avss.n76 10.4659
R638 avss.n256 avss.n255 10.4659
R639 avss.n186 avss.n79 10.4659
R640 avss.n187 avss.n100 10.4659
R641 avss.n238 avss.n237 10.4659
R642 avss.n211 avss.n103 10.4659
R643 avss.n150 avss.n131 10.4659
R644 avss.n166 avss.n165 10.4659
R645 avss.n169 avss.n168 10.4659
R646 avss.n173 avss.n119 10.4659
R647 avss.n193 avss.n192 10.4659
R648 avss.n196 avss.n195 10.4659
R649 avss.n199 avss.n198 10.4659
R650 avss.n206 avss.n205 10.4659
R651 avss.n212 avss.n24 10.4574
R652 avss.n329 avss.n328 10.4488
R653 avss.n333 avss.n20 10.4301
R654 avss.n201 avss.n26 10.4152
R655 avss.n335 avss.n334 10.3988
R656 avss.n226 avss.n225 10.3825
R657 avss.n113 avss.n108 10.3825
R658 avss.n244 avss.n243 10.3825
R659 avss.n184 avss.n86 10.3825
R660 avss.n125 avss.n84 10.3825
R661 avss.n262 avss.n261 10.3825
R662 avss.n142 avss.n63 10.3825
R663 avss.n336 avss.n13 10.3029
R664 avss.n233 avss.n232 10.3029
R665 avss.n242 avss.n96 10.3029
R666 avss.n245 avss.n90 10.3029
R667 avss.n251 avss.n250 10.3029
R668 avss.n260 avss.n72 10.3029
R669 avss.n263 avss.n66 10.3029
R670 avss.n285 avss.n284 10.3029
R671 avss.n60 avss.n53 9.81158
R672 avss.n171 avss.n89 9.70903
R673 avss.t69 avss.t98 9.61512
R674 avss.n171 avss.n65 9.37433
R675 avss.n298 avss.t112 6.99295
R676 avss.n128 avss.t66 6.99295
R677 avss.n268 avss.n267 6.53477
R678 avss.n201 avss.n20 6.4005
R679 avss.n336 avss.n335 6.32245
R680 avss.n232 avss.n226 6.32245
R681 avss.n113 avss.n96 6.32245
R682 avss.n245 avss.n244 6.32245
R683 avss.n250 avss.n86 6.32245
R684 avss.n125 avss.n72 6.32245
R685 avss.n263 avss.n262 6.32245
R686 avss.n284 avss.n63 6.32245
R687 avss.n341 avss.n11 6.29691
R688 avss.n287 avss.n60 4.94826
R689 avss.n306 avss.n305 3.79309
R690 avss.n320 avss.n29 3.5246
R691 avss.n37 avss.n29 3.5246
R692 avss.n30 avss.n28 3.5246
R693 avss.n37 avss.n28 3.5246
R694 avss.n4 avss.n2 3.5246
R695 avss.n154 avss.n4 3.5246
R696 avss.n267 avss.n3 3.5246
R697 avss.n154 avss.n3 3.5246
R698 avss.n271 avss.n270 3.07647
R699 avss.n350 avss.n349 2.90959
R700 avss.n173 avss.n172 2.6571
R701 avss.n64 avss.n60 2.3284
R702 avss.n344 avss.n343 2.3255
R703 avss.n47 avss.n46 2.3255
R704 avss.n303 avss.n34 2.3255
R705 avss.n278 avss.n277 2.24027
R706 avss.n10 avss 2.08383
R707 avss.n275 avss.n273 2.05988
R708 avss.n278 avss.n276 2.05939
R709 avss.n307 avss.n47 1.38845
R710 avss.n274 avss.n273 1.25531
R711 avss.n337 avss.n336 1.163
R712 avss.n232 avss.n231 1.163
R713 avss.n227 avss.n96 1.163
R714 avss.n246 avss.n245 1.163
R715 avss.n250 avss.n249 1.163
R716 avss.n87 avss.n72 1.163
R717 avss.n264 avss.n263 1.163
R718 avss.n284 avss.n283 1.163
R719 avss.n20 avss.n19 1.163
R720 avss.n343 avss.n342 1.1255
R721 avss.n305 avss.n32 1.03383
R722 avss.n304 avss.n303 0.925801
R723 avss.n282 avss.n64 0.606932
R724 avss.n229 avss.n1 0.577925
R725 avss.n268 avss.n266 0.577925
R726 avss.n19 avss.n9 0.563
R727 avss.n228 avss.n227 0.563
R728 avss.n231 avss.n230 0.563
R729 avss.n338 avss.n337 0.563
R730 avss.n88 avss.n87 0.563
R731 avss.n249 avss.n248 0.563
R732 avss.n247 avss.n246 0.563
R733 avss.n283 avss.n282 0.563
R734 avss.n265 avss.n264 0.563
R735 avss.n351 avss.n350 0.494944
R736 avss.n272 avss.n271 0.494944
R737 avss.n319 avss.n318 0.4655
R738 avss.n340 avss.n339 0.401201
R739 avss.n281 avss.n272 0.356756
R740 avss.n340 avss.n0 0.304064
R741 avss.n287 avss.n286 0.287571
R742 avss.n342 avss.n9 0.243877
R743 avss.n248 avss.n88 0.230632
R744 avss.n248 avss.n247 0.230632
R745 avss.n247 avss.n89 0.204142
R746 avss.n279 avss.n278 0.181204
R747 avss.n294 avss.n53 0.163374
R748 avss.n280 avss.n12 0.163113
R749 avss.n172 avss.n171 0.143769
R750 avss.n341 avss.n340 0.128227
R751 avss.n313 avss.n41 0.119019
R752 avss avss.n351 0.106457
R753 avss.n88 avss.n65 0.104391
R754 avss.n12 avss.n0 0.0954724
R755 avss.n11 avss.n10 0.068442
R756 avss.n281 avss.n280 0.058173
R757 avss.n46 avss.n32 0.048994
R758 avss.n230 avss.n228 0.0444317
R759 avss.n266 avss.n265 0.0418243
R760 avss.n339 avss.n338 0.0386637
R761 avss.n10 avss 0.0334815
R762 avss.n317 avss.n34 0.0319759
R763 avss.t86 avss.n274 0.0307671
R764 avss.n339 avss.n9 0.0307152
R765 avss.n338 avss.n12 0.0278388
R766 avss.n265 avss.n65 0.0245992
R767 avss.t6 avss.n275 0.0217969
R768 avss.t89 avss.n276 0.0217969
R769 avss.n277 avss.t75 0.0217969
R770 avss.n280 avss.n279 0.0211667
R771 avss.n275 avss.t86 0.0183453
R772 avss.n276 avss.t6 0.0183453
R773 avss.n277 avss.t89 0.0183453
R774 avss.n230 avss.n229 0.0170139
R775 avss.n34 avss.n33 0.0164639
R776 avss.n318 avss.n32 0.0161626
R777 avss.n342 avss.n341 0.0108477
R778 avss.n274 avss.t149 0.0103017
R779 avss.n33 avss.n11 0.0068253
R780 avss.n228 avss.n89 0.00555689
R781 avss.n272 avss 0.00344634
R782 avss.n282 avss.n281 0.00302845
R783 avss.n279 avss.n273 0.000669675
R784 avss.n318 avss.n317 0.000650602
R785 avss.n351 avss.n0 0.000606383
R786 avss.n229 avss.n12 0.000579014
R787 avss.n281 avss.n266 0.000579014
R788 ena.n5 ena.t2 396.2
R789 ena.n5 ena.t3 381.825
R790 ena.n1 ena.t5 305.348
R791 ena.n0 ena.t6 302.945
R792 ena.n3 ena.t4 196.596
R793 ena.n2 ena.t0 112.272
R794 ena.n2 ena.t1 110.207
R795 ena.n5 ena.n4 4.5005
R796 ena.n4 ena.n3 2.03668
R797 ena.n4 ena.n1 1.72267
R798 ena.n3 ena.n2 1.20571
R799 ena.n1 ena.n0 1.06763
R800 ena.n0 ena 0.368556
R801 ena ena.n5 0.062375
R802 a_3638_4788.t1 a_3638_4788.t3 660.754
R803 a_3638_4788.t3 a_3638_4788.t0 235.388
R804 a_3638_4788.t3 a_3638_4788.t4 107.769
R805 a_3638_4788.t3 a_3638_4788.t2 105.281
R806 a_4194_4788.t0 a_4194_4788.t4 660.745
R807 a_4194_4788.t4 a_4194_4788.t1 235.613
R808 a_4194_4788.t4 a_4194_4788.t2 107.96
R809 a_4194_4788.t4 a_4194_4788.t3 105.281
R810 a_2368_4788.n1 a_2368_4788.t2 660.24
R811 a_2368_4788.t1 a_2368_4788.n1 660.24
R812 a_2368_4788.n1 a_2368_4788.t3 236.429
R813 a_2368_4788.n0 a_2368_4788.t9 107.941
R814 a_2368_4788.n1 a_2368_4788.t0 106.373
R815 a_2368_4788.n0 a_2368_4788.t7 106.373
R816 a_2368_4788.n0 a_2368_4788.t6 106.373
R817 a_2368_4788.n0 a_2368_4788.t8 106.373
R818 a_2368_4788.n0 a_2368_4788.t4 106.373
R819 a_2368_4788.n0 a_2368_4788.t5 106.373
R820 a_2368_4788.n0 a_2368_4788.t10 106.373
R821 a_2368_4788.n1 a_2368_4788.n0 11.6107
R822 avdd.n245 avdd.n244 32453.4
R823 avdd.n244 avdd.n230 32453.4
R824 avdd.n246 avdd.n245 22625.9
R825 avdd.n298 avdd.n230 22623
R826 avdd.n243 avdd.n228 17294.1
R827 avdd.n243 avdd.n240 17294.1
R828 avdd.n247 avdd.n240 12162.6
R829 avdd.n299 avdd.n228 12161
R830 avdd.n298 avdd.n297 8083.85
R831 avdd.n246 avdd.n231 8069.1
R832 avdd.n297 avdd.n296 6124.84
R833 avdd.n299 avdd.n229 4569.24
R834 avdd.n248 avdd.n247 4561.54
R835 avdd.n248 avdd.n232 3771.24
R836 avdd.n232 avdd.n229 3765.08
R837 avdd.n296 avdd.n231 3546.27
R838 avdd.n242 avdd.n241 1252.21
R839 avdd.n226 avdd.n0 1014.54
R840 avdd.n241 avdd.n239 949.297
R841 avdd.n154 avdd.n144 841.241
R842 avdd.n154 avdd.n145 841.241
R843 avdd.n144 avdd.n143 841.241
R844 avdd.n145 avdd.n143 841.241
R845 avdd.n172 avdd.n120 841.241
R846 avdd.n172 avdd.n121 841.241
R847 avdd.n171 avdd.n121 841.241
R848 avdd.n171 avdd.n120 841.241
R849 avdd.n177 avdd.n114 841.241
R850 avdd.n177 avdd.n115 841.241
R851 avdd.n115 avdd.n113 841.241
R852 avdd.n114 avdd.n113 841.241
R853 avdd.n196 avdd.n87 841.241
R854 avdd.n185 avdd.n87 841.241
R855 avdd.n185 avdd.n88 841.241
R856 avdd.n196 avdd.n88 841.241
R857 avdd.n201 avdd.n83 841.241
R858 avdd.n199 avdd.n83 841.241
R859 avdd.n200 avdd.n199 841.241
R860 avdd.n201 avdd.n200 841.241
R861 avdd.n211 avdd.n21 841.241
R862 avdd.n211 avdd.n22 841.241
R863 avdd.n210 avdd.n22 841.241
R864 avdd.n210 avdd.n21 841.241
R865 avdd.n216 avdd.n17 841.241
R866 avdd.n216 avdd.n18 841.241
R867 avdd.n18 avdd.n11 841.241
R868 avdd.n17 avdd.n11 841.241
R869 avdd.n141 avdd.n139 841.241
R870 avdd.n155 avdd.n139 841.241
R871 avdd.n155 avdd.n138 841.241
R872 avdd.n141 avdd.n138 841.241
R873 avdd.n128 avdd.n123 841.241
R874 avdd.n128 avdd.n124 841.241
R875 avdd.n134 avdd.n124 841.241
R876 avdd.n134 avdd.n123 841.241
R877 avdd.n110 avdd.n109 841.241
R878 avdd.n178 avdd.n110 841.241
R879 avdd.n179 avdd.n178 841.241
R880 avdd.n179 avdd.n109 841.241
R881 avdd.n187 avdd.n99 841.241
R882 avdd.n188 avdd.n187 841.241
R883 avdd.n188 avdd.n86 841.241
R884 avdd.n99 avdd.n86 841.241
R885 avdd.n85 avdd.n81 841.241
R886 avdd.n85 avdd.n82 841.241
R887 avdd.n203 avdd.n82 841.241
R888 avdd.n203 avdd.n81 841.241
R889 avdd.n28 avdd.n24 841.241
R890 avdd.n28 avdd.n25 841.241
R891 avdd.n32 avdd.n25 841.241
R892 avdd.n32 avdd.n24 841.241
R893 avdd.n217 avdd.n13 841.241
R894 avdd.n15 avdd.n13 841.241
R895 avdd.n15 avdd.n12 841.241
R896 avdd.n217 avdd.n12 841.241
R897 avdd.n56 avdd.n49 841.241
R898 avdd.n53 avdd.n49 841.241
R899 avdd.n56 avdd.n48 841.241
R900 avdd.n70 avdd.n43 841.241
R901 avdd.n70 avdd.n44 841.241
R902 avdd.n43 avdd.n42 841.241
R903 avdd.n44 avdd.n42 841.241
R904 avdd.n40 avdd.n37 841.241
R905 avdd.n40 avdd.n38 841.241
R906 avdd.n71 avdd.n38 841.241
R907 avdd.n71 avdd.n37 841.241
R908 avdd.n266 avdd.n264 841.241
R909 avdd.n275 avdd.n264 841.241
R910 avdd.n275 avdd.n269 841.241
R911 avdd.n269 avdd.n266 841.241
R912 avdd.n285 avdd.n256 841.241
R913 avdd.n286 avdd.n256 841.241
R914 avdd.n285 avdd.n257 841.241
R915 avdd.n286 avdd.n257 841.241
R916 avdd.n272 avdd.n234 841.241
R917 avdd.n272 avdd.n235 841.241
R918 avdd.n294 avdd.n235 841.241
R919 avdd.n294 avdd.n234 841.241
R920 avdd.n277 avdd.n259 841.241
R921 avdd.n281 avdd.n259 841.241
R922 avdd.n277 avdd.n260 841.241
R923 avdd.n281 avdd.n260 841.241
R924 avdd.n301 avdd.n226 757.859
R925 avdd.n167 avdd.t18 660.576
R926 avdd.n167 avdd.t16 660.562
R927 avdd.n5 avdd.t4 660.562
R928 avdd.n94 avdd.t6 660.562
R929 avdd.n106 avdd.t10 660.562
R930 avdd.n165 avdd.t8 660.562
R931 avdd.n221 avdd.t12 660.562
R932 avdd.n4 avdd.t2 660.562
R933 avdd.n206 avdd.t14 660.562
R934 avdd.n253 avdd.t20 660.391
R935 avdd.n290 avdd.t22 660.38
R936 avdd.n249 avdd.n239 338.13
R937 avdd.n55 avdd.n39 311.062
R938 avdd.n300 avdd.n227 305.512
R939 avdd.n250 avdd.n249 230.186
R940 avdd.n251 avdd.n238 179.423
R941 avdd.n296 avdd.n295 168.218
R942 avdd.t23 avdd.n55 149.226
R943 avdd.t3 avdd.n39 149.226
R944 avdd.t3 avdd.n41 149.226
R945 avdd.t1 avdd.n14 149.226
R946 avdd.t1 avdd.n16 149.226
R947 avdd.t11 avdd.n23 149.226
R948 avdd.t11 avdd.n26 149.226
R949 avdd.n202 avdd.t13 149.226
R950 avdd.n198 avdd.t13 149.226
R951 avdd.n197 avdd.t5 149.226
R952 avdd.n186 avdd.t5 149.226
R953 avdd.t9 avdd.n101 149.226
R954 avdd.t9 avdd.n112 149.226
R955 avdd.t7 avdd.n122 149.226
R956 avdd.t7 avdd.n125 149.226
R957 avdd.t15 avdd.n140 149.226
R958 avdd.t15 avdd.n142 149.226
R959 avdd.n54 avdd.n48 145.906
R960 avdd.n41 avdd.n14 133.113
R961 avdd.n23 avdd.n16 133.113
R962 avdd.n202 avdd.n26 133.113
R963 avdd.n198 avdd.n197 133.113
R964 avdd.n186 avdd.n101 133.113
R965 avdd.n122 avdd.n112 133.113
R966 avdd.n140 avdd.n125 133.113
R967 avdd.t17 avdd.n258 128.886
R968 avdd.t17 avdd.n261 128.886
R969 avdd.t19 avdd.n233 125.255
R970 avdd.n273 avdd.t21 125.255
R971 avdd.n147 avdd.n137 114.112
R972 avdd.n152 avdd.n147 112.749
R973 avdd.n274 avdd.n258 111.338
R974 avdd.n135 avdd.n126 91.9447
R975 avdd.n181 avdd.n180 91.9447
R976 avdd.n97 avdd.n95 91.9447
R977 avdd.n33 avdd.n7 91.9447
R978 avdd.n34 avdd.n10 91.9447
R979 avdd.n62 avdd.n61 91.9447
R980 avdd.n136 avdd.n131 91.9447
R981 avdd.n205 avdd.n204 91.9447
R982 avdd.n207 avdd.n30 90.0623
R983 avdd.n164 avdd.n118 90.0623
R984 avdd.n182 avdd.n105 90.0623
R985 avdd.n195 avdd.n194 90.0623
R986 avdd.n220 avdd.n6 90.0623
R987 avdd.n65 avdd.n64 90.0623
R988 avdd.n60 avdd.n59 90.0623
R989 avdd.n168 avdd.n130 90.0623
R990 avdd.n169 avdd.n129 85.4593
R991 avdd.n163 avdd.n162 85.4593
R992 avdd.n183 avdd.n100 85.4593
R993 avdd.n193 avdd.n192 85.4593
R994 avdd.n208 avdd.n29 85.4593
R995 avdd.n219 avdd.n9 85.4593
R996 avdd.n58 avdd.n46 85.4593
R997 avdd.n66 avdd.n35 85.4593
R998 avdd.n158 avdd.n129 85.0829
R999 avdd.n160 avdd.n135 85.0829
R1000 avdd.n162 avdd.n161 85.0829
R1001 avdd.n180 avdd.n108 85.0829
R1002 avdd.n100 avdd.n98 85.0829
R1003 avdd.n190 avdd.n97 85.0829
R1004 avdd.n192 avdd.n191 85.0829
R1005 avdd.n79 avdd.n29 85.0829
R1006 avdd.n77 avdd.n33 85.0829
R1007 avdd.n74 avdd.n34 85.0829
R1008 avdd.n76 avdd.n9 85.0829
R1009 avdd.n51 avdd.n46 85.0829
R1010 avdd.n73 avdd.n35 85.0829
R1011 avdd.n61 avdd.n36 85.0829
R1012 avdd.n157 avdd.n136 85.0829
R1013 avdd.n204 avdd.n80 85.0829
R1014 avdd.n169 avdd.n127 83.9534
R1015 avdd.n163 avdd.n117 83.9534
R1016 avdd.n184 avdd.n183 83.9534
R1017 avdd.n193 avdd.n84 83.9534
R1018 avdd.n208 avdd.n27 83.9534
R1019 avdd.n219 avdd.n8 83.9534
R1020 avdd.n67 avdd.n66 83.9534
R1021 avdd.n89 avdd.n30 82.824
R1022 avdd.n127 avdd.n119 82.824
R1023 avdd.n174 avdd.n118 82.824
R1024 avdd.n175 avdd.n117 82.824
R1025 avdd.n116 avdd.n105 82.824
R1026 avdd.n184 avdd.n103 82.824
R1027 avdd.n195 avdd.n93 82.824
R1028 avdd.n92 avdd.n84 82.824
R1029 avdd.n27 avdd.n20 82.824
R1030 avdd.n213 avdd.n6 82.824
R1031 avdd.n64 avdd.n19 82.824
R1032 avdd.n214 avdd.n8 82.824
R1033 avdd.n68 avdd.n67 82.824
R1034 avdd.n59 avdd.n45 82.824
R1035 avdd.n146 avdd.n130 82.824
R1036 avdd.n47 avdd.n45 64.4732
R1037 avdd.n265 avdd.n263 51.1301
R1038 avdd.n282 avdd.n280 50.4217
R1039 avdd.n242 avdd.n0 49.7553
R1040 avdd.n57 avdd.n56 46.2505
R1041 avdd.n56 avdd.t23 46.2505
R1042 avdd.n218 avdd.n217 46.2505
R1043 avdd.n217 avdd.t1 46.2505
R1044 avdd.n209 avdd.n24 46.2505
R1045 avdd.t11 avdd.n24 46.2505
R1046 avdd.n81 avdd.n31 46.2505
R1047 avdd.t13 avdd.n81 46.2505
R1048 avdd.n104 avdd.n99 46.2505
R1049 avdd.n99 avdd.t5 46.2505
R1050 avdd.n109 avdd.n107 46.2505
R1051 avdd.t9 avdd.n109 46.2505
R1052 avdd.n170 avdd.n123 46.2505
R1053 avdd.t7 avdd.n123 46.2505
R1054 avdd.n149 avdd.n141 46.2505
R1055 avdd.t15 avdd.n141 46.2505
R1056 avdd.n218 avdd.n11 46.2505
R1057 avdd.t1 avdd.n11 46.2505
R1058 avdd.n210 avdd.n209 46.2505
R1059 avdd.t11 avdd.n210 46.2505
R1060 avdd.n200 avdd.n31 46.2505
R1061 avdd.n200 avdd.t13 46.2505
R1062 avdd.n104 avdd.n88 46.2505
R1063 avdd.n88 avdd.t5 46.2505
R1064 avdd.n113 avdd.n107 46.2505
R1065 avdd.t9 avdd.n113 46.2505
R1066 avdd.n171 avdd.n170 46.2505
R1067 avdd.t7 avdd.n171 46.2505
R1068 avdd.n149 avdd.n143 46.2505
R1069 avdd.t15 avdd.n143 46.2505
R1070 avdd.n63 avdd.n42 46.2505
R1071 avdd.t3 avdd.n42 46.2505
R1072 avdd.n63 avdd.n40 46.2505
R1073 avdd.t3 avdd.n40 46.2505
R1074 avdd.n70 avdd.n69 46.2505
R1075 avdd.t3 avdd.n70 46.2505
R1076 avdd.n216 avdd.n215 46.2505
R1077 avdd.t1 avdd.n216 46.2505
R1078 avdd.n212 avdd.n211 46.2505
R1079 avdd.n211 avdd.t11 46.2505
R1080 avdd.n91 avdd.n83 46.2505
R1081 avdd.n83 avdd.t13 46.2505
R1082 avdd.n102 avdd.n87 46.2505
R1083 avdd.n87 avdd.t5 46.2505
R1084 avdd.n177 avdd.n176 46.2505
R1085 avdd.t9 avdd.n177 46.2505
R1086 avdd.n173 avdd.n172 46.2505
R1087 avdd.n172 avdd.t7 46.2505
R1088 avdd.n154 avdd.n153 46.2505
R1089 avdd.t15 avdd.n154 46.2505
R1090 avdd.n53 avdd.n52 46.2505
R1091 avdd.n72 avdd.n71 46.2505
R1092 avdd.n71 avdd.t3 46.2505
R1093 avdd.n75 avdd.n15 46.2505
R1094 avdd.t1 avdd.n15 46.2505
R1095 avdd.n78 avdd.n25 46.2505
R1096 avdd.t11 avdd.n25 46.2505
R1097 avdd.n96 avdd.n82 46.2505
R1098 avdd.t13 avdd.n82 46.2505
R1099 avdd.n189 avdd.n188 46.2505
R1100 avdd.n188 avdd.t5 46.2505
R1101 avdd.n178 avdd.n111 46.2505
R1102 avdd.n178 avdd.t9 46.2505
R1103 avdd.n159 avdd.n124 46.2505
R1104 avdd.t7 avdd.n124 46.2505
R1105 avdd.n156 avdd.n155 46.2505
R1106 avdd.n155 avdd.t15 46.2505
R1107 avdd.n267 avdd.n234 46.2505
R1108 avdd.t19 avdd.n234 46.2505
R1109 avdd.n237 avdd.n235 46.2505
R1110 avdd.t19 avdd.n235 46.2505
R1111 avdd.n287 avdd.n286 46.2505
R1112 avdd.n286 avdd.t17 46.2505
R1113 avdd.n269 avdd.n268 46.2505
R1114 avdd.t21 avdd.n269 46.2505
R1115 avdd.n280 avdd.n259 46.2505
R1116 avdd.t17 avdd.n259 46.2505
R1117 avdd.n264 avdd.n263 46.2505
R1118 avdd.t21 avdd.n264 46.2505
R1119 avdd.n285 avdd.n284 46.2505
R1120 avdd.t17 avdd.n285 46.2505
R1121 avdd.n284 avdd.n260 46.2505
R1122 avdd.t17 avdd.n260 46.2505
R1123 avdd.n52 avdd.n50 44.9285
R1124 avdd.n156 avdd.n137 39.8981
R1125 avdd.n50 avdd.n47 39.5797
R1126 avdd.n153 avdd.n152 39.2634
R1127 avdd.n50 avdd.n48 37.0005
R1128 avdd.n49 avdd.n46 37.0005
R1129 avdd.n55 avdd.n49 37.0005
R1130 avdd.n34 avdd.n12 37.0005
R1131 avdd.n14 avdd.n12 37.0005
R1132 avdd.n13 avdd.n9 37.0005
R1133 avdd.n16 avdd.n13 37.0005
R1134 avdd.n33 avdd.n32 37.0005
R1135 avdd.n32 avdd.n23 37.0005
R1136 avdd.n29 avdd.n28 37.0005
R1137 avdd.n28 avdd.n26 37.0005
R1138 avdd.n192 avdd.n85 37.0005
R1139 avdd.n198 avdd.n85 37.0005
R1140 avdd.n97 avdd.n86 37.0005
R1141 avdd.n197 avdd.n86 37.0005
R1142 avdd.n187 avdd.n100 37.0005
R1143 avdd.n187 avdd.n186 37.0005
R1144 avdd.n180 avdd.n179 37.0005
R1145 avdd.n179 avdd.n101 37.0005
R1146 avdd.n162 avdd.n110 37.0005
R1147 avdd.n112 avdd.n110 37.0005
R1148 avdd.n135 avdd.n134 37.0005
R1149 avdd.n134 avdd.n122 37.0005
R1150 avdd.n129 avdd.n128 37.0005
R1151 avdd.n128 avdd.n125 37.0005
R1152 avdd.n148 avdd.n139 37.0005
R1153 avdd.n142 avdd.n139 37.0005
R1154 avdd.n64 avdd.n17 37.0005
R1155 avdd.n17 avdd.n14 37.0005
R1156 avdd.n18 avdd.n8 37.0005
R1157 avdd.n18 avdd.n16 37.0005
R1158 avdd.n21 avdd.n6 37.0005
R1159 avdd.n23 avdd.n21 37.0005
R1160 avdd.n27 avdd.n22 37.0005
R1161 avdd.n26 avdd.n22 37.0005
R1162 avdd.n201 avdd.n30 37.0005
R1163 avdd.n202 avdd.n201 37.0005
R1164 avdd.n199 avdd.n84 37.0005
R1165 avdd.n199 avdd.n198 37.0005
R1166 avdd.n196 avdd.n195 37.0005
R1167 avdd.n197 avdd.n196 37.0005
R1168 avdd.n185 avdd.n184 37.0005
R1169 avdd.n186 avdd.n185 37.0005
R1170 avdd.n114 avdd.n105 37.0005
R1171 avdd.n114 avdd.n101 37.0005
R1172 avdd.n117 avdd.n115 37.0005
R1173 avdd.n115 avdd.n112 37.0005
R1174 avdd.n120 avdd.n118 37.0005
R1175 avdd.n122 avdd.n120 37.0005
R1176 avdd.n127 avdd.n121 37.0005
R1177 avdd.n125 avdd.n121 37.0005
R1178 avdd.n151 avdd.n145 37.0005
R1179 avdd.n145 avdd.n142 37.0005
R1180 avdd.n67 avdd.n44 37.0005
R1181 avdd.n44 avdd.n41 37.0005
R1182 avdd.n38 avdd.n35 37.0005
R1183 avdd.n41 avdd.n38 37.0005
R1184 avdd.n61 avdd.n37 37.0005
R1185 avdd.n39 avdd.n37 37.0005
R1186 avdd.n59 avdd.n43 37.0005
R1187 avdd.n43 avdd.n39 37.0005
R1188 avdd.n144 avdd.n130 37.0005
R1189 avdd.n144 avdd.n140 37.0005
R1190 avdd.n138 avdd.n136 37.0005
R1191 avdd.n140 avdd.n138 37.0005
R1192 avdd.n204 avdd.n203 37.0005
R1193 avdd.n203 avdd.n202 37.0005
R1194 avdd.n294 avdd.n293 37.0005
R1195 avdd.n295 avdd.n294 37.0005
R1196 avdd.n266 avdd.n265 37.0005
R1197 avdd.n266 avdd.n233 37.0005
R1198 avdd.n282 avdd.n281 37.0005
R1199 avdd.n281 avdd.n261 37.0005
R1200 avdd.n276 avdd.n275 37.0005
R1201 avdd.n275 avdd.n274 37.0005
R1202 avdd.n278 avdd.n277 37.0005
R1203 avdd.n277 avdd.n258 37.0005
R1204 avdd.n272 avdd.n271 37.0005
R1205 avdd.n273 avdd.n272 37.0005
R1206 avdd.n271 avdd.n256 37.0005
R1207 avdd.n258 avdd.n256 37.0005
R1208 avdd.n257 avdd.n254 37.0005
R1209 avdd.n261 avdd.n257 37.0005
R1210 avdd.n54 avdd.n53 36.2372
R1211 avdd.n51 avdd.n36 35.7439
R1212 avdd.n296 avdd.n232 35.604
R1213 avdd.n288 avdd.n287 26.6196
R1214 avdd.n292 avdd.n237 25.9151
R1215 avdd.n238 avdd.n227 25.2054
R1216 avdd.n60 avdd.n58 24.1639
R1217 avdd.n150 avdd.n148 24.0137
R1218 avdd.n151 avdd.n150 23.5906
R1219 avdd.n280 avdd.n279 23.2301
R1220 avdd.n279 avdd.n263 23.2301
R1221 avdd.n293 avdd.n236 23.1206
R1222 avdd.n293 avdd.n292 23.0608
R1223 avdd.n283 avdd.n282 23.0608
R1224 avdd.n283 avdd.n254 23.0608
R1225 avdd.n265 avdd.n236 22.7005
R1226 avdd.n288 avdd.n254 21.9434
R1227 avdd.n287 avdd.n255 20.2328
R1228 avdd.n255 avdd.n237 20.2328
R1229 avdd.n271 avdd.n262 19.0862
R1230 avdd.n69 avdd.n45 17.1477
R1231 avdd.n69 avdd.n68 17.1477
R1232 avdd.n215 avdd.n19 17.1477
R1233 avdd.n215 avdd.n214 17.1477
R1234 avdd.n213 avdd.n212 17.1477
R1235 avdd.n212 avdd.n20 17.1477
R1236 avdd.n92 avdd.n91 17.1477
R1237 avdd.n102 avdd.n93 17.1477
R1238 avdd.n103 avdd.n102 17.1477
R1239 avdd.n176 avdd.n116 17.1477
R1240 avdd.n176 avdd.n175 17.1477
R1241 avdd.n174 avdd.n173 17.1477
R1242 avdd.n173 avdd.n119 17.1477
R1243 avdd.n153 avdd.n146 17.1477
R1244 avdd.n52 avdd.n51 17.1477
R1245 avdd.n72 avdd.n36 17.1477
R1246 avdd.n73 avdd.n72 17.1477
R1247 avdd.n75 avdd.n74 17.1477
R1248 avdd.n76 avdd.n75 17.1477
R1249 avdd.n78 avdd.n77 17.1477
R1250 avdd.n79 avdd.n78 17.1477
R1251 avdd.n96 avdd.n80 17.1477
R1252 avdd.n191 avdd.n96 17.1477
R1253 avdd.n190 avdd.n189 17.1477
R1254 avdd.n189 avdd.n98 17.1477
R1255 avdd.n111 avdd.n108 17.1477
R1256 avdd.n161 avdd.n111 17.1477
R1257 avdd.n160 avdd.n159 17.1477
R1258 avdd.n159 avdd.n158 17.1477
R1259 avdd.n157 avdd.n156 17.1477
R1260 avdd.n279 avdd.n278 16.2647
R1261 avdd.n68 avdd.n19 15.2961
R1262 avdd.n214 avdd.n213 15.2961
R1263 avdd.n89 avdd.n20 15.2961
R1264 avdd.n93 avdd.n92 15.2961
R1265 avdd.n116 avdd.n103 15.2961
R1266 avdd.n175 avdd.n174 15.2961
R1267 avdd.n146 avdd.n119 15.2961
R1268 avdd.n74 avdd.n73 15.2961
R1269 avdd.n77 avdd.n76 15.2961
R1270 avdd.n80 avdd.n79 15.2961
R1271 avdd.n191 avdd.n190 15.2961
R1272 avdd.n108 avdd.n98 15.2961
R1273 avdd.n161 avdd.n160 15.2961
R1274 avdd.n158 avdd.n157 15.2961
R1275 avdd.n267 avdd.n236 15.193
R1276 avdd.n284 avdd.n283 14.8746
R1277 avdd.n150 avdd.n149 14.4286
R1278 avdd.n276 avdd.n262 13.2702
R1279 avdd.n170 avdd.n169 11.9584
R1280 avdd.n163 avdd.n107 11.9584
R1281 avdd.n183 avdd.n104 11.9584
R1282 avdd.n193 avdd.n31 11.9584
R1283 avdd.n209 avdd.n208 11.9584
R1284 avdd.n219 avdd.n218 11.9584
R1285 avdd.n66 avdd.n63 11.9584
R1286 avdd.n58 avdd.n57 11.9302
R1287 avdd.n284 avdd.n262 11.6153
R1288 avdd.n268 avdd.n262 11.365
R1289 avdd.n90 avdd.n89 10.8684
R1290 avdd.n169 avdd.n168 9.77806
R1291 avdd.n164 avdd.n163 9.77806
R1292 avdd.n183 avdd.n182 9.77806
R1293 avdd.n194 avdd.n193 9.77806
R1294 avdd.n208 avdd.n207 9.77806
R1295 avdd.n220 avdd.n219 9.77806
R1296 avdd.n66 avdd.n65 9.77806
R1297 avdd.n271 avdd.n270 8.8005
R1298 avdd.n148 avdd.n137 8.25174
R1299 avdd.n152 avdd.n151 8.14595
R1300 avdd.t23 avdd.n54 8.02261
R1301 avdd.n270 avdd.n255 7.6005
R1302 avdd.n91 avdd.n90 6.27974
R1303 avdd.n249 avdd.n248 6.16717
R1304 avdd.n248 avdd.n231 6.16717
R1305 avdd.n229 avdd.n227 6.16717
R1306 avdd.n297 avdd.n229 6.16717
R1307 avdd.n250 avdd.n232 4.74409
R1308 avdd.n295 avdd.n233 3.63107
R1309 avdd.t21 avdd.t19 3.63107
R1310 avdd.n274 avdd.n273 3.63107
R1311 avdd.n150 avdd.n147 3.36892
R1312 avdd.n247 avdd.n239 3.36414
R1313 avdd.n247 avdd.n246 3.36414
R1314 avdd.n300 avdd.n299 3.36414
R1315 avdd.n299 avdd.n298 3.36414
R1316 avdd.n289 avdd.n288 3.10844
R1317 avdd.n292 avdd.n291 3.1005
R1318 avdd.n251 avdd.n250 2.57768
R1319 avdd.n57 avdd.n47 2.51578
R1320 avdd.n252 avdd.n225 1.34749
R1321 avdd.n243 avdd.n242 1.20965
R1322 avdd.n244 avdd.n243 1.20965
R1323 avdd.n306 avdd.n0 1.13445
R1324 avdd.n241 avdd.n240 1.05164
R1325 avdd.n245 avdd.n240 1.05164
R1326 avdd.n228 avdd.n226 1.05164
R1327 avdd.n230 avdd.n228 1.05164
R1328 avdd.n270 avdd.n253 0.9305
R1329 avdd.n291 avdd.n252 0.877364
R1330 avdd.n165 avdd.n164 0.7755
R1331 avdd.n182 avdd.n106 0.7755
R1332 avdd.n194 avdd.n94 0.7755
R1333 avdd.n221 avdd.n220 0.7755
R1334 avdd.n65 avdd.n4 0.7755
R1335 avdd.n60 avdd.n5 0.7755
R1336 avdd.n168 avdd.n167 0.7755
R1337 avdd.n207 avdd.n206 0.7755
R1338 avdd.n301 avdd.n300 0.621859
R1339 avdd.n2 avdd.n1 0.552286
R1340 avdd.n238 avdd.n225 0.504
R1341 avdd.n302 avdd.n301 0.490106
R1342 avdd.n206 avdd.n3 0.3755
R1343 avdd.n132 avdd.n94 0.3755
R1344 avdd.n166 avdd.n106 0.3755
R1345 avdd.n166 avdd.n165 0.3755
R1346 avdd.n167 avdd.n166 0.3755
R1347 avdd.n222 avdd.n5 0.3755
R1348 avdd.n222 avdd.n4 0.3755
R1349 avdd.n222 avdd.n221 0.3755
R1350 avdd.n268 avdd.n267 0.359379
R1351 avdd.n149 avdd.n131 0.281202
R1352 avdd.n170 avdd.n126 0.281202
R1353 avdd.n181 avdd.n107 0.281202
R1354 avdd.n104 avdd.n95 0.281202
R1355 avdd.n205 avdd.n31 0.281202
R1356 avdd.n209 avdd.n7 0.281202
R1357 avdd.n218 avdd.n10 0.281202
R1358 avdd.n63 avdd.n62 0.281202
R1359 avdd.n304 avdd.n303 0.27802
R1360 avdd.n303 avdd.n225 0.244654
R1361 avdd.n132 avdd.n3 0.244171
R1362 avdd.n252 avdd.n251 0.233
R1363 avdd.n224 avdd.n2 0.221333
R1364 avdd.n306 avdd.n305 0.192137
R1365 avdd.n305 avdd.n304 0.185806
R1366 avdd.n90 avdd.n2 0.172219
R1367 avdd.n133 avdd.n132 0.14963
R1368 avdd.n291 avdd.n290 0.122295
R1369 avdd.n223 avdd.n3 0.121149
R1370 avdd.n290 avdd.n289 0.119303
R1371 avdd.n278 avdd.n276 0.117931
R1372 avdd.n303 avdd.n302 0.090332
R1373 avdd.n305 avdd.n1 0.0714439
R1374 avdd.n304 avdd.n224 0.0714439
R1375 avdd.n164 avdd.n126 0.0573889
R1376 avdd.n182 avdd.n181 0.0573889
R1377 avdd.n194 avdd.n95 0.0573889
R1378 avdd.n220 avdd.n7 0.0573889
R1379 avdd.n65 avdd.n10 0.0573889
R1380 avdd.n62 avdd.n60 0.0573889
R1381 avdd.n168 avdd.n131 0.0573889
R1382 avdd.n207 avdd.n205 0.0573889
R1383 avdd.n133 avdd.n1 0.0547069
R1384 avdd.n224 avdd.n223 0.0547069
R1385 avdd avdd.n306 0.0146048
R1386 avdd.n289 avdd 0.0139615
R1387 avdd.n290 avdd.n253 0.00377715
R1388 avdd.n302 avdd 0.00325827
R1389 avdd.n166 avdd.n133 0.000801568
R1390 avdd.n223 avdd.n222 0.000801568
R1391 level_shifter_0.outb_h.n0 level_shifter_0.outb_h.t1 660.24
R1392 level_shifter_0.outb_h.n0 level_shifter_0.outb_h.t0 235.004
R1393 level_shifter_0.outb_h level_shifter_0.outb_h.t2 127.82
R1394 level_shifter_0.outb_h.n0 level_shifter_0.outb_h.t3 116.334
R1395 level_shifter_0.outb_h.n0 level_shifter_0.outb_h.t4 107.222
R1396 level_shifter_0.outb_h level_shifter_0.outb_h.n0 11.5134
R1397 level_shifter_0.out_h level_shifter_0.out_h.t0 660.24
R1398 level_shifter_0.out_h level_shifter_0.out_h.t1 235.251
R1399 level_shifter_0.out_h level_shifter_0.out_h.t4 116.338
R1400 level_shifter_0.out_h.n0 level_shifter_0.out_h.t2 110.648
R1401 level_shifter_0.out_h level_shifter_0.out_h.t5 106.773
R1402 level_shifter_0.out_h.n0 level_shifter_0.out_h.t6 106.382
R1403 level_shifter_0.out_h.n0 level_shifter_0.out_h.t3 104.746
R1404 level_shifter_0.out_h level_shifter_0.out_h.n0 21.9372
R1405 a_3082_4788.t0 a_3082_4788.t2 660.769
R1406 a_3082_4788.t2 a_3082_4788.t1 235.127
R1407 a_3082_4788.t2 a_3082_4788.t3 107.582
R1408 a_3082_4788.t2 a_3082_4788.t4 105.273
R1409 dvdd.n18 dvdd.n13 1312.94
R1410 dvdd.n22 dvdd.n12 1312.94
R1411 dvdd.n22 dvdd.n13 1312.94
R1412 dvdd.n5 dvdd.n4 1312.94
R1413 dvdd.n26 dvdd.n25 1108.24
R1414 dvdd.n25 dvdd.n8 1108.24
R1415 dvdd.n6 dvdd.n5 704.168
R1416 dvdd.n34 dvdd.n3 697.11
R1417 dvdd.n37 dvdd.t6 668.082
R1418 dvdd.n0 dvdd.t3 662.312
R1419 dvdd.n31 dvdd.n3 596.572
R1420 dvdd.n31 dvdd.n6 589.715
R1421 dvdd.n26 dvdd.n6 497.647
R1422 dvdd.n8 dvdd.n3 497.647
R1423 dvdd.n24 dvdd.n23 345.777
R1424 dvdd.n32 dvdd.t2 334.182
R1425 dvdd.n24 dvdd.t2 332.08
R1426 dvdd.t4 dvdd.n32 332.08
R1427 dvdd.n33 dvdd.n4 277.072
R1428 dvdd.n23 dvdd.t0 264.262
R1429 dvdd.n18 dvdd.n17 237.584
R1430 dvdd.n39 dvdd.t5 228.498
R1431 dvdd.n9 dvdd.t1 228.239
R1432 dvdd.n20 dvdd.n19 137.024
R1433 dvdd.t4 dvdd.n5 106.007
R1434 dvdd.n19 dvdd.n16 100.001
R1435 dvdd.n20 dvdd.n12 95.2318
R1436 dvdd.n16 dvdd.n13 92.5005
R1437 dvdd.n13 dvdd.t0 92.5005
R1438 dvdd.n27 dvdd.n26 92.5005
R1439 dvdd.n26 dvdd.t2 92.5005
R1440 dvdd.n35 dvdd.n34 92.5005
R1441 dvdd.n28 dvdd.n5 92.5005
R1442 dvdd.n14 dvdd.n8 92.5005
R1443 dvdd.n8 dvdd.t2 92.5005
R1444 dvdd.n28 dvdd.n2 90.9905
R1445 dvdd.n29 dvdd.n28 75.1118
R1446 dvdd.n34 dvdd.n33 74.3381
R1447 dvdd.n17 dvdd.n12 70.7763
R1448 dvdd.n30 dvdd.n29 62.9034
R1449 dvdd.n25 dvdd.n11 61.6672
R1450 dvdd.n25 dvdd.n24 61.6672
R1451 dvdd.n30 dvdd.n1 57.4176
R1452 dvdd.n27 dvdd.n7 53.0829
R1453 dvdd.n29 dvdd.n27 53.0829
R1454 dvdd.n35 dvdd.n2 52.7584
R1455 dvdd.n19 dvdd.n18 46.2505
R1456 dvdd.n4 dvdd.n2 46.2505
R1457 dvdd.n31 dvdd.n30 46.2505
R1458 dvdd.n32 dvdd.n31 46.2505
R1459 dvdd.n22 dvdd.n21 46.2505
R1460 dvdd.n23 dvdd.n22 46.2505
R1461 dvdd.n21 dvdd.n20 44.1706
R1462 dvdd.n15 dvdd.n14 40.0601
R1463 dvdd.n16 dvdd.n15 23.8938
R1464 dvdd.n33 dvdd.t4 21.4216
R1465 dvdd.n17 dvdd.t0 16.7394
R1466 dvdd.n36 dvdd.n1 13.4634
R1467 dvdd.n14 dvdd.n1 12.4864
R1468 dvdd.n11 dvdd.n10 9.51845
R1469 dvdd.n15 dvdd.n11 3.41383
R1470 dvdd.n37 dvdd.n36 2.3255
R1471 dvdd.n10 dvdd.n7 1.83845
R1472 dvdd.n10 dvdd.n9 1.55446
R1473 dvdd.n21 dvdd.n7 0.459987
R1474 dvdd.n39 dvdd.n38 0.317167
R1475 dvdd.n40 dvdd.n39 0.153726
R1476 dvdd.n40 dvdd.n0 0.146137
R1477 dvdd.n36 dvdd.n35 0.129793
R1478 dvdd.n9 dvdd.n0 0.0618011
R1479 dvdd.n38 dvdd.n37 0.038
R1480 dvdd.n41 dvdd.n40 0.0228214
R1481 dvdd dvdd.n41 0.0228214
R1482 dvdd.n38 dvdd 0.004875
R1483 dvdd.n41 dvdd 0.001125
R1484 a_4750_4788.t1 a_4750_4788.t2 660.756
R1485 a_4750_4788.t2 a_4750_4788.t0 235.773
R1486 a_4750_4788.t2 a_4750_4788.t3 108.153
R1487 a_4750_4788.t2 a_4750_4788.t4 105.281
R1488 a_1414_4786.n0 a_1414_4786.t2 237.433
R1489 a_1414_4786.n0 a_1414_4786.t3 235.407
R1490 a_1414_4786.t1 a_1414_4786.n0 233.657
R1491 a_1414_4786.n0 a_1414_4786.t10 113.971
R1492 a_1414_4786.n0 a_1414_4786.t4 105.537
R1493 a_1414_4786.n0 a_1414_4786.t0 104.177
R1494 a_1414_4786.n0 a_1414_4786.t6 104.175
R1495 a_1414_4786.n0 a_1414_4786.t5 104.175
R1496 a_1414_4786.n0 a_1414_4786.t8 104.175
R1497 a_1414_4786.n0 a_1414_4786.t11 104.175
R1498 a_1414_4786.n0 a_1414_4786.t7 104.175
R1499 a_1414_4786.n0 a_1414_4786.t9 104.175
R1500 a_5306_4788.t1 a_5306_4788.t2 660.806
R1501 a_5306_4788.t2 a_5306_4788.t0 235.982
R1502 a_5306_4788.t2 a_5306_4788.t3 108.346
R1503 a_5306_4788.t2 a_5306_4788.t4 105.281
R1504 dvss.n42 dvss.n38 25476.2
R1505 dvss.n43 dvss.n19 9928.12
R1506 dvss.n62 dvss.n11 2126.44
R1507 dvss.n24 dvss.n11 2126.44
R1508 dvss.n62 dvss.n12 2126.44
R1509 dvss.n24 dvss.n12 2126.44
R1510 dvss.n40 dvss.n35 1836.74
R1511 dvss.n44 dvss.n35 1836.74
R1512 dvss.n44 dvss.n34 1836.74
R1513 dvss.n37 dvss.n9 1836.74
R1514 dvss.n65 dvss.n9 1836.74
R1515 dvss.n37 dvss.n10 1836.74
R1516 dvss.n65 dvss.n10 1836.74
R1517 dvss.n54 dvss.n22 1790.38
R1518 dvss.n22 dvss.n20 1790.38
R1519 dvss.n21 dvss.n20 1790.38
R1520 dvss.n54 dvss.n21 1790.38
R1521 dvss.n64 dvss.n63 1740.52
R1522 dvss.n25 dvss.n23 1449.84
R1523 dvss.n56 dvss.n17 1407.97
R1524 dvss.n56 dvss.n18 1407.97
R1525 dvss.n49 dvss.n17 1407.97
R1526 dvss.n49 dvss.n18 1407.97
R1527 dvss.t2 dvss.n43 818.846
R1528 dvss.n41 dvss.n40 776.158
R1529 dvss.n38 dvss.t0 667.819
R1530 dvss.n64 dvss.t0 667.819
R1531 dvss.n27 dvss.n26 592.715
R1532 dvss.n63 dvss.t4 569.837
R1533 dvss.n48 dvss.t3 468.853
R1534 dvss.n55 dvss.t6 367.87
R1535 dvss.n42 dvss.n41 329.875
R1536 dvss.n26 dvss.t4 317.377
R1537 dvss.n41 dvss.n34 316.318
R1538 dvss.n13 dvss.n11 294.214
R1539 dvss.n10 dvss.n8 292.5
R1540 dvss.t0 dvss.n10 292.5
R1541 dvss.n9 dvss.n7 292.5
R1542 dvss.t0 dvss.n9 292.5
R1543 dvss.n40 dvss.n39 292.5
R1544 dvss.n45 dvss.n44 292.5
R1545 dvss.n44 dvss.t2 292.5
R1546 dvss.n18 dvss.n15 292.5
R1547 dvss.t3 dvss.n18 292.5
R1548 dvss.n54 dvss.n53 292.5
R1549 dvss.t6 dvss.n54 292.5
R1550 dvss.n50 dvss.n49 292.5
R1551 dvss.n49 dvss.n48 292.5
R1552 dvss.n31 dvss.n17 292.5
R1553 dvss.t3 dvss.n17 292.5
R1554 dvss.n30 dvss.n20 292.5
R1555 dvss.t6 dvss.n20 292.5
R1556 dvss.n57 dvss.n56 292.5
R1557 dvss.n56 dvss.n55 292.5
R1558 dvss.n60 dvss.n12 292.5
R1559 dvss.n12 dvss.t4 292.5
R1560 dvss.n11 dvss.t4 292.5
R1561 dvss.n26 dvss.n25 252.459
R1562 dvss.n6 dvss.t7 239.136
R1563 dvss.t2 dvss.n42 233.216
R1564 dvss.n1 dvss.t1 229.315
R1565 dvss.n34 dvss.n33 195.184
R1566 dvss.n66 dvss.n65 195
R1567 dvss.n65 dvss.n64 195
R1568 dvss.n37 dvss.n36 195
R1569 dvss.n38 dvss.n37 195
R1570 dvss.n35 dvss.n32 195
R1571 dvss.n43 dvss.n35 195
R1572 dvss.n52 dvss.n22 195
R1573 dvss.n48 dvss.n22 195
R1574 dvss.n28 dvss.n21 195
R1575 dvss.n23 dvss.n21 195
R1576 dvss.n23 dvss.n19 155.083
R1577 dvss.n24 dvss.n14 146.25
R1578 dvss.n25 dvss.n24 146.25
R1579 dvss.n62 dvss.n61 146.25
R1580 dvss.n63 dvss.n62 146.25
R1581 dvss.n61 dvss.n60 138.166
R1582 dvss.n53 dvss.n52 116.504
R1583 dvss.t6 dvss.t3 100.984
R1584 dvss.n47 dvss.n46 97.6305
R1585 dvss.n61 dvss.n13 86.5887
R1586 dvss.n36 dvss.n8 86.1306
R1587 dvss.n3 dvss.t5 84.1047
R1588 dvss.n39 dvss.n33 81.8974
R1589 dvss.n36 dvss.n7 74.9169
R1590 dvss.n45 dvss.n33 74.0493
R1591 dvss.n52 dvss.n51 57.0188
R1592 dvss.n58 dvss.n57 55.3148
R1593 dvss.n53 dvss.n29 53.0829
R1594 dvss.n60 dvss.n59 53.0829
R1595 dvss.n50 dvss.n47 48.155
R1596 dvss.n55 dvss.n19 46.8857
R1597 dvss.n39 dvss.n32 43.9756
R1598 dvss.n51 dvss.n50 42.7064
R1599 dvss.n66 dvss.n8 39.1038
R1600 dvss.n30 dvss.n16 31.8699
R1601 dvss.n57 dvss.n16 26.2862
R1602 dvss.n68 dvss.n67 17.1865
R1603 dvss.n46 dvss.n45 17.0668
R1604 dvss.n29 dvss.n6 14.0183
R1605 dvss.n68 dvss.n7 13.3694
R1606 dvss.n46 dvss.n32 12.1441
R1607 dvss.n27 dvss.n16 11.3033
R1608 dvss.n59 dvss.n58 10.109
R1609 dvss.n51 dvss.n31 6.79342
R1610 dvss.n59 dvss.n14 6.606
R1611 dvss.n5 dvss.n0 5.813
R1612 dvss.n58 dvss.n15 5.62852
R1613 dvss.n13 dvss.n2 5.6005
R1614 dvss.n29 dvss.n28 4.75646
R1615 dvss.n67 dvss.n1 4.6505
R1616 dvss.n67 dvss.n66 2.95435
R1617 dvss.n3 dvss.n0 2.6255
R1618 dvss.n70 dvss.n2 2.33934
R1619 dvss.n27 dvss.n2 1.88621
R1620 dvss.n69 dvss.n68 1.82171
R1621 dvss.n31 dvss.n30 1.46336
R1622 dvss.n69 dvss.n6 1.44933
R1623 dvss.n4 dvss.n3 1.2505
R1624 dvss.n47 dvss.n15 1.09622
R1625 dvss.n5 dvss 0.8755
R1626 dvss.n4 dvss 0.583833
R1627 dvss.n72 dvss.n0 0.438
R1628 dvss.n28 dvss.n27 0.26472
R1629 dvss.n69 dvss 0.119327
R1630 dvss.n70 dvss.n69 0.0769887
R1631 dvss.n16 dvss.n14 0.0592156
R1632 dvss.n71 dvss.n1 0.0536915
R1633 dvss.n70 dvss.n5 0.0472557
R1634 dvss.n71 dvss.n70 0.0133337
R1635 dvss.n72 dvss.n71 0.0125637
R1636 dvss.n5 dvss.n4 0.0019313
R1637 dvss dvss.n72 0.00178337
R1638 dvss.n4 dvss 0.000977099
R1639 dout.n1 dout.t2 243.876
R1640 dout.n0 dout.t1 230.631
R1641 dout.n0 dout.t0 228.215
R1642 dout.n1 dout.n0 3.11789
R1643 dout dout.n1 0.306432
R1644 a_2982_4700.t1 a_2982_4700.n0 661.461
R1645 a_2982_4700.n0 a_2982_4700.t0 236.12
R1646 a_2982_4700.n0 a_2982_4700.t3 108.308
R1647 a_2982_4700.n0 a_2982_4700.t5 107.8
R1648 a_2982_4700.n1 a_2982_4700.t2 107.362
R1649 a_2982_4700.n1 a_2982_4700.t4 105.01
R1650 a_2982_4700.n0 a_2982_4700.n1 16.7414
C0 a_6490_9768# a_6158_9768# 0.307869f
C1 level_shifter_0.out_h a_2526_4188# 0.106807f
C2 avss a_7984_7168# 0.209517f
C3 avdd a_9664_3118# 0.031575f
C4 a_11636_7168# a_10660_3118# 0.018676f
C5 avdd a_6086_5653# 0.788381f
C6 avdd a_6178_518# 0.012005f
C7 dout dvdd 0.892013f
C8 a_6988_7168# a_6656_7168# 0.307869f
C9 a_11324_3118# ena 2.91e-19
C10 avss a_11304_7168# 0.145925f
C11 a_5348_3118# a_5016_3118# 0.307869f
C12 a_4830_9768# avss 0.142763f
C13 a_10474_9768# a_10142_9768# 0.307869f
C14 dout ena 0.18382f
C15 a_9830_518# a_9498_518# 0.307869f
C16 avdd level_shifter_0.out_h 2.25409f
C17 level_shifter_0.inb_l a_8714_4659# 0.012649f
C18 avdd a_1510_9768# 0.071412f
C19 avss a_4020_3118# 0.365534f
C20 avdd a_6510_518# 0.012005f
C21 a_3006_5653# a_3622_5653# 0.00665f
C22 avss a_9482_5327# 0.007616f
C23 avss a_10308_7168# 0.144844f
C24 avss a_9332_3118# 0.214403f
C25 a_4592_4788# level_shifter_0.out_h 0.001601f
C26 avdd a_3522_518# 0.012005f
C27 avdd a_4850_518# 0.012005f
C28 a_1178_9768# avdd 0.071412f
C29 avdd a_3004_7168# 0.548273f
C30 a_11636_7168# a_11304_7168# 0.307345f
C31 level_shifter_0.outb_h a_7560_4786# 0.017545f
C32 a_7718_4786# avdd 0.60786f
C33 avss a_9664_3118# 0.211499f
C34 a_6178_518# avss 0.184675f
C35 avss a_6086_5653# 0.001818f
C36 a_1862_518# a_1530_518# 0.307869f
C37 a_10162_518# a_9830_518# 0.307869f
C38 avdd a_7818_9768# 0.071412f
C39 avss level_shifter_0.out_h 4.25651f
C40 avss a_1510_9768# 0.142763f
C41 a_6510_518# avss 0.184675f
C42 a_7340_3118# a_7008_3118# 0.307869f
C43 level_shifter_0.outb_h a_1364_3118# 1.01e-19
C44 avdd a_5494_9768# 0.071412f
C45 avss a_3522_518# 0.184675f
C46 avdd a_8980_7168# 0.049449f
C47 a_10640_7168# a_10308_7168# 0.307869f
C48 a_8502_518# a_8834_518# 0.307869f
C49 a_5470_5653# a_4854_5653# 0.00665f
C50 avss a_4850_518# 0.184675f
C51 a_7154_9768# a_6822_9768# 0.307869f
C52 a_1178_9768# avss 0.142763f
C53 a_3004_7168# avss 0.209517f
C54 level_shifter_0.outb_h a_3480_4788# 0.018927f
C55 a_7718_4786# avss 0.630608f
C56 a_10826_518# a_10494_518# 0.307869f
C57 a_11636_7168# level_shifter_0.out_h 3.09e-21
C58 avdd a_8336_3118# 0.032475f
C59 avdd a_1198_518# 0.012005f
C60 avdd a_10142_9768# 0.071412f
C61 a_9996_3118# a_9664_3118# 0.307869f
C62 a_4664_7168# a_4332_7168# 0.307869f
C63 a_7818_9768# avss 0.142763f
C64 a_6324_7168# a_6656_7168# 0.307869f
C65 a_9644_7168# a_9312_7168# 0.307869f
C66 avss a_6260_4788# 0.892467f
C67 avss a_5494_9768# 0.142763f
C68 a_7718_4786# a_11636_7168# 0.04522f
C69 level_shifter_0.outb_h a_8004_3118# 1.78e-19
C70 avdd a_4000_7168# 0.385508f
C71 a_4036_4788# a_3480_4788# 0.009712f
C72 avss a_8980_7168# 0.243852f
C73 avdd a_2174_9768# 0.071412f
C74 a_3006_5653# level_shifter_0.out_h 2.23e-19
C75 a_2028_3118# a_1696_3118# 0.307869f
C76 a_8336_3118# avss 0.220223f
C77 a_1198_518# avss 0.184675f
C78 a_11890_5939# dvdd 0.120615f
C79 dvdd a_7984_7168# 0.001364f
C80 avdd a_9498_518# 0.012005f
C81 avss a_10142_9768# 0.142763f
C82 a_11890_5939# ena 0.177772f
C83 avss a_7672_3118# 0.28253f
C84 avdd a_7838_518# 0.012005f
C85 level_shifter_0.outb_h a_5148_4788# 0.018927f
C86 a_10806_9768# a_10474_9768# 0.307869f
C87 avdd a_11490_518# 0.031753f
C88 a_8668_3118# a_9000_3118# 0.307869f
C89 a_10992_3118# avdd 0.009316f
C90 avss a_4000_7168# 0.209517f
C91 a_9482_5327# ena 0.117123f
C92 avss a_2174_9768# 0.142763f
C93 a_4830_9768# a_4498_9768# 0.307869f
C94 avdd level_shifter_0.inb_l 0.368358f
C95 avdd a_10162_518# 0.012005f
C96 a_6490_9768# a_6822_9768# 0.307869f
C97 avss a_9498_518# 0.184675f
C98 level_shifter_0.outb_h a_4036_4788# 0.018927f
C99 a_9810_9768# a_9478_9768# 0.307869f
C100 a_5862_4788# a_7560_4786# 3.04e-20
C101 a_9664_3118# ena 1.38e-20
C102 a_11158_518# a_11490_518# 0.307869f
C103 avss a_7838_518# 0.184675f
C104 dvdd level_shifter_0.out_h 0.040401f
C105 avdd a_5992_7168# 0.548273f
C106 avss a_11490_518# 0.348069f
C107 ena level_shifter_0.out_h 0.3516f
C108 level_shifter_0.out_h a_2924_4788# 0.001827f
C109 a_10992_3118# avss 0.20921f
C110 a_11890_5939# dout 0.638473f
C111 a_5846_518# a_5514_518# 0.307869f
C112 level_shifter_0.inb_l avss 0.875565f
C113 a_3854_518# a_3522_518# 0.307869f
C114 dout a_11304_7168# 7.41e-20
C115 a_3668_7168# a_3336_7168# 0.307869f
C116 a_10162_518# avss 0.184675f
C117 a_5470_5653# a_6086_5653# 0.00665f
C118 a_7718_4786# dvdd 1.2174f
C119 avdd a_8170_518# 0.012005f
C120 a_7718_4786# ena 0.523822f
C121 level_shifter_0.outb_h a_8714_4659# 0.229072f
C122 avdd a_7506_518# 0.012005f
C123 a_10992_3118# a_11636_7168# 0.018676f
C124 avdd a_10806_9768# 0.071412f
C125 a_1178_9768# a_846_9768# 0.307869f
C126 avss a_5992_7168# 0.209517f
C127 avss a_1696_3118# 0.533397f
C128 level_shifter_0.inb_l a_11636_7168# 0.164792f
C129 avdd a_7486_9768# 0.071412f
C130 a_6260_4788# ena 5.02e-21
C131 avdd a_6988_7168# 0.342919f
C132 a_8648_7168# a_8980_7168# 0.307869f
C133 a_514_7168# a_680_7168# 0.311537f
C134 dout level_shifter_0.out_h 6.46e-21
C135 a_8170_518# avss 0.184675f
C136 avdd a_4332_7168# 0.070399f
C137 avdd a_9000_3118# 0.032475f
C138 avss a_7506_518# 0.184675f
C139 a_6676_3118# avss 0.739782f
C140 avss a_10806_9768# 0.142763f
C141 avdd a_7560_4786# 0.026816f
C142 a_7672_3118# ena 1.82e-19
C143 a_9644_7168# a_9976_7168# 0.307869f
C144 avdd a_2506_9768# 0.071412f
C145 a_5862_4788# level_shifter_0.outb_h 0.140134f
C146 avss a_7486_9768# 0.142763f
C147 avdd a_10972_7168# 0.609955f
C148 a_3834_9768# a_3502_9768# 0.307869f
C149 a_6012_3118# a_5680_3118# 0.307869f
C150 a_7718_4786# dout 1.09434f
C151 a_2858_518# a_3190_518# 0.307869f
C152 a_4020_3118# a_3688_3118# 0.307869f
C153 a_1032_3118# a_1364_3118# 0.307869f
C154 avss a_6988_7168# 0.209517f
C155 a_2194_518# a_1862_518# 0.307869f
C156 avdd a_8502_518# 0.012005f
C157 avdd a_5846_518# 0.012005f
C158 avss a_4332_7168# 0.209517f
C159 avss a_9000_3118# 0.215061f
C160 a_10162_518# a_10494_518# 0.307869f
C161 a_7506_518# a_7174_518# 0.307869f
C162 a_3004_7168# a_3336_7168# 0.307869f
C163 avdd a_8814_9768# 0.071412f
C164 avss a_7560_4786# 0.445517f
C165 a_9498_518# a_9166_518# 0.307869f
C166 a_8814_9768# a_9146_9768# 0.307869f
C167 avdd a_9644_7168# 0.305891f
C168 avss a_2506_9768# 0.142763f
C169 avdd a_1530_518# 0.012005f
C170 avss a_10972_7168# 0.144844f
C171 a_5704_4788# level_shifter_0.out_h 0.001092f
C172 avdd a_1862_518# 0.012005f
C173 a_6510_518# a_6842_518# 0.307869f
C174 a_8502_518# avss 0.184675f
C175 a_10992_3118# ena 2.52e-20
C176 a_1364_3118# avss 0.282494f
C177 level_shifter_0.inb_l dvdd 0.663728f
C178 level_shifter_0.inb_l a_8648_7168# 3.07e-19
C179 avdd a_6324_7168# 0.548273f
C180 avdd a_4238_5653# 0.701946f
C181 avss a_5846_518# 0.184675f
C182 level_shifter_0.inb_l ena 1.01705f
C183 avss a_8814_9768# 0.142763f
C184 a_9810_9768# a_10142_9768# 0.307869f
C185 a_6988_7168# a_7320_7168# 0.307869f
C186 avdd a_514_9768# 0.091264f
C187 avss a_3480_4788# 0.828006f
C188 level_shifter_0.outb_h a_2526_4188# 0.017016f
C189 avdd a_2672_7168# 0.548273f
C190 a_514_7168# level_shifter_0.out_h 0.142627f
C191 avss a_9644_7168# 0.198487f
C192 a_3024_3118# a_3356_3118# 0.307869f
C193 avdd a_3190_518# 0.012005f
C194 avss a_1530_518# 0.184675f
C195 avdd a_6656_7168# 0.548273f
C196 a_2360_3118# a_2028_3118# 0.307869f
C197 avss a_1862_518# 0.184675f
C198 avdd level_shifter_0.outb_h 1.603f
C199 avdd a_10328_3118# 0.009597f
C200 a_3170_9768# a_3502_9768# 0.307869f
C201 a_10640_7168# a_10972_7168# 0.307869f
C202 a_5704_4788# a_6260_4788# 0.009712f
C203 avss a_6324_7168# 0.209517f
C204 a_7672_3118# a_7340_3118# 0.307869f
C205 avss a_4238_5653# 0.00413f
C206 level_shifter_0.outb_h a_4592_4788# 0.018927f
C207 a_5148_4788# a_4592_4788# 0.009712f
C208 a_4518_518# a_4186_518# 0.307869f
C209 avdd a_8834_518# 0.012005f
C210 avss a_8004_3118# 0.241301f
C211 a_1012_7168# a_1344_7168# 0.307869f
C212 avdd a_9312_7168# 0.056717f
C213 a_5862_4788# a_6702_5653# 0.11184f
C214 a_9664_3118# a_9332_3118# 0.307869f
C215 a_514_9768# avss 0.305402f
C216 a_10992_3118# a_11324_3118# 0.307869f
C217 avdd a_3502_9768# 0.071412f
C218 avss a_2672_7168# 0.209517f
C219 avdd a_1842_9768# 0.071412f
C220 a_5182_518# a_5514_518# 0.307869f
C221 avdd a_8316_7168# 0.04813f
C222 a_9482_5327# level_shifter_0.out_h 0.102468f
C223 a_7718_4786# a_11890_5939# 0.052047f
C224 avss a_3190_518# 0.184675f
C225 avss a_6656_7168# 0.209517f
C226 level_shifter_0.inb_l dout 0.13931f
C227 a_6676_3118# a_7008_3118# 0.307869f
C228 level_shifter_0.outb_h avss 4.51566f
C229 a_10328_3118# avss 0.20921f
C230 avss a_5148_4788# 0.865328f
C231 a_4036_4788# a_4592_4788# 0.009712f
C232 avss a_5680_3118# 0.739782f
C233 a_7154_9768# a_7486_9768# 0.307869f
C234 avss a_8834_518# 0.184675f
C235 a_7718_4786# a_9482_5327# 1.23e-19
C236 a_6178_518# a_6510_518# 0.307869f
C237 avss a_9312_7168# 0.243852f
C238 a_3024_3118# avss 0.739899f
C239 avdd a_4664_7168# 0.061398f
C240 avss a_3502_9768# 0.142763f
C241 avss a_1842_9768# 0.142763f
C242 avdd a_4518_518# 0.012005f
C243 avss a_8316_7168# 0.243852f
C244 level_shifter_0.outb_h a_11636_7168# 7.58e-20
C245 a_10806_9768# a_11138_9768# 0.307869f
C246 a_11636_7168# a_10328_3118# 0.00554f
C247 avss a_4036_4788# 0.823951f
C248 a_7560_4786# ena 0.161553f
C249 avdd a_8714_4659# 0.401456f
C250 avss a_4352_3118# 0.350904f
C251 a_10972_7168# ena 6.11e-20
C252 a_1178_9768# a_1510_9768# 0.307869f
C253 a_7718_4786# level_shifter_0.out_h 0.144107f
C254 a_4684_3118# a_4352_3118# 0.307869f
C255 a_10328_3118# a_9996_3118# 0.307869f
C256 a_2526_518# a_2858_518# 0.307869f
C257 a_4000_7168# a_3668_7168# 0.307869f
C258 avdd a_5162_9768# 0.071412f
C259 avdd a_5826_9768# 0.071412f
C260 avss a_2360_3118# 0.739899f
C261 a_5348_3118# a_5680_3118# 0.307869f
C262 a_4664_7168# avss 0.209517f
C263 level_shifter_0.outb_h a_3006_5653# 9.7e-22
C264 avdd a_6702_5653# 0.791907f
C265 a_4518_518# avss 0.184675f
C266 avdd a_9830_518# 0.012005f
C267 avdd a_1344_7168# 0.049439f
C268 avdd a_3834_9768# 0.071412f
C269 a_6260_4788# level_shifter_0.out_h 9.06e-20
C270 a_9644_7168# dvdd 4.86e-19
C271 a_2924_4788# a_3480_4788# 0.009712f
C272 avss a_8714_4659# 0.033517f
C273 a_9644_7168# ena 1.74e-20
C274 a_10992_3118# a_10660_3118# 0.307869f
C275 avdd a_8668_3118# 0.032475f
C276 avdd a_8150_9768# 0.071412f
C277 a_5182_518# avdd 0.012005f
C278 a_866_518# avdd 0.012005f
C279 a_2672_7168# a_2340_7168# 0.307869f
C280 avdd a_5514_518# 0.012005f
C281 a_1012_7168# avdd 0.050125f
C282 avdd a_11470_9768# 0.090673f
C283 a_2526_518# a_2194_518# 0.307869f
C284 a_6344_3118# a_6676_3118# 0.307869f
C285 a_5862_4788# avdd 0.82569f
C286 avss a_5162_9768# 0.142763f
C287 avss a_5826_9768# 0.142763f
C288 avdd a_2858_518# 0.012005f
C289 avdd a_10474_9768# 0.071412f
C290 a_8004_3118# ena 0.010181f
C291 avdd a_7652_7168# 0.056845f
C292 avss a_6702_5653# 0.001818f
C293 avss a_9830_518# 0.184675f
C294 avss a_1344_7168# 0.239502f
C295 avss a_3834_9768# 0.142763f
C296 level_shifter_0.inb_l a_11890_5939# 9.85e-21
C297 a_5660_7168# a_5992_7168# 0.307869f
C298 avdd a_5328_7168# 0.436049f
C299 a_8668_3118# avss 0.217285f
C300 a_4166_9768# a_3834_9768# 0.307869f
C301 avss a_8150_9768# 0.142763f
C302 a_5182_518# avss 0.184675f
C303 a_514_9768# a_846_9768# 0.307869f
C304 a_2692_3118# a_3024_3118# 0.307869f
C305 level_shifter_0.outb_h dvdd 0.015582f
C306 a_866_518# avss 0.184675f
C307 avdd a_2526_518# 0.012005f
C308 avdd a_4186_518# 0.012005f
C309 avss a_5514_518# 0.184675f
C310 a_1012_7168# avss 0.239502f
C311 avss a_6012_3118# 0.739782f
C312 level_shifter_0.outb_h ena 0.463304f
C313 avss a_11470_9768# 0.307678f
C314 level_shifter_0.outb_h a_2924_4788# 0.018927f
C315 a_5862_4788# avss 1.04054f
C316 level_shifter_0.inb_l a_9482_5327# 4.08e-19
C317 level_shifter_0.inb_l a_10308_7168# 1.8e-19
C318 avdd a_9976_7168# 0.609955f
C319 a_2858_518# avss 0.184675f
C320 avdd a_2194_518# 0.012005f
C321 avss a_10474_9768# 0.142763f
C322 a_7652_7168# avss 0.209517f
C323 a_9312_7168# ena 3.61e-19
C324 a_9166_518# a_8834_518# 0.307869f
C325 a_8648_7168# a_8316_7168# 0.307869f
C326 a_2838_9768# a_2506_9768# 0.307869f
C327 avss a_2028_3118# 0.739899f
C328 avss a_5328_7168# 0.209517f
C329 avdd a_3170_9768# 0.071412f
C330 a_2692_3118# a_2360_3118# 0.307869f
C331 level_shifter_0.inb_l level_shifter_0.out_h 0.255743f
C332 avss a_4186_518# 0.184675f
C333 a_2526_518# avss 0.184675f
C334 avdd a_2008_7168# 0.066489f
C335 avss a_9976_7168# 0.144844f
C336 a_5826_9768# a_6158_9768# 0.307869f
C337 avss a_2194_518# 0.184675f
C338 avss a_3356_3118# 0.66303f
C339 level_shifter_0.outb_h dout 1.42e-20
C340 a_7718_4786# level_shifter_0.inb_l 0.881308f
C341 avdd a_9146_9768# 0.071412f
C342 a_4238_5653# a_4854_5653# 0.00665f
C343 a_3170_9768# avss 0.142763f
C344 a_1032_3118# a_700_3118# 0.307869f
C345 avss a_2526_4188# 0.699047f
C346 avdd a_700_3118# 0.308767f
C347 a_8714_4659# ena 0.035705f
C348 a_7652_7168# a_7320_7168# 0.307869f
C349 avss a_2008_7168# 0.209517f
C350 avdd a_11158_518# 0.012005f
C351 a_1032_3118# avss 0.614509f
C352 avdd avss 0.348303p
C353 a_8814_9768# a_8482_9768# 0.307869f
C354 a_9332_3118# a_9000_3118# 0.307869f
C355 avss a_4592_4788# 0.824116f
C356 avdd a_4166_9768# 0.071412f
C357 dvdd a_6702_5653# 0.004947f
C358 a_10972_7168# a_11304_7168# 0.307869f
C359 avss a_9146_9768# 0.142763f
C360 a_3622_5653# a_4238_5653# 0.00665f
C361 avss a_700_3118# 0.725885f
C362 avdd a_11636_7168# 1.3903f
C363 avss a_11158_518# 0.184675f
C364 a_5862_4788# dvdd 0.00524f
C365 avdd a_7174_518# 0.012005f
C366 level_shifter_0.outb_h a_5704_4788# 0.018927f
C367 a_5148_4788# a_5704_4788# 0.009712f
C368 a_5862_4788# ena 0.002113f
C369 a_4684_3118# avss 0.334568f
C370 avdd a_9996_3118# 0.015329f
C371 a_7560_4786# level_shifter_0.out_h 0.001495f
C372 avss a_4166_9768# 0.142763f
C373 avdd a_10640_7168# 0.609955f
C374 a_7818_9768# a_7486_9768# 0.307869f
C375 avdd a_7320_7168# 0.065995f
C376 a_6178_518# a_5846_518# 0.307869f
C377 avdd a_3006_5653# 0.816596f
C378 a_11636_7168# avss 0.808235f
C379 level_shifter_0.outb_h a_514_7168# 0.068229f
C380 a_10328_3118# a_10660_3118# 0.307869f
C381 a_7718_4786# a_7560_4786# 0.015996f
C382 a_4186_518# a_3854_518# 0.307869f
C383 avss a_7174_518# 0.184675f
C384 a_11138_9768# a_11470_9768# 0.307869f
C385 avdd a_6158_9768# 0.071412f
C386 level_shifter_0.out_h a_3480_4788# 0.001602f
C387 avss a_9996_3118# 0.20921f
C388 avdd a_10494_518# 0.012005f
C389 avss a_10640_7168# 0.144844f
C390 a_2008_7168# a_2340_7168# 0.307869f
C391 a_5348_3118# avss 0.693821f
C392 avdd a_2340_7168# 0.399783f
C393 avss a_7320_7168# 0.209517f
C394 a_1676_7168# a_1344_7168# 0.307869f
C395 a_3006_5653# avss 0.002318f
C396 level_shifter_0.outb_h a_9482_5327# 0.202516f
C397 level_shifter_0.outb_h a_9332_3118# 3.26e-19
C398 a_8170_518# a_7838_518# 0.307869f
C399 a_2924_4788# a_2526_4188# 0.031652f
C400 a_7718_4786# a_9644_7168# 2.34e-20
C401 a_8316_7168# a_7984_7168# 0.307869f
C402 a_7506_518# a_7838_518# 0.307869f
C403 a_866_518# a_534_518# 0.307869f
C404 avss a_6158_9768# 0.142763f
C405 avdd dvdd 1.48803f
C406 avdd a_8648_7168# 0.047906f
C407 avss a_10494_518# 0.184675f
C408 a_4664_7168# a_4996_7168# 0.307869f
C409 a_4000_7168# a_4332_7168# 0.307869f
C410 avdd a_3854_518# 0.012005f
C411 avdd a_2924_4788# 0.003752f
C412 avdd ena 1.6305f
C413 avdd a_7154_9768# 0.071412f
C414 avdd a_9166_518# 0.012005f
C415 avss a_2340_7168# 0.209517f
C416 a_6344_3118# a_6012_3118# 0.307869f
C417 level_shifter_0.outb_h level_shifter_0.out_h 3.79716f
C418 avdd a_846_9768# 0.071412f
C419 a_2692_3118# avss 0.739899f
C420 a_5148_4788# level_shifter_0.out_h 0.001601f
C421 avdd a_4498_9768# 0.071412f
C422 a_4352_3118# a_4020_3118# 0.307869f
C423 a_3522_518# a_3190_518# 0.307869f
C424 a_3004_7168# a_2672_7168# 0.307869f
C425 avdd a_5470_5653# 0.761298f
C426 a_2174_9768# a_2506_9768# 0.307869f
C427 avss a_8648_7168# 0.243852f
C428 avss dvdd 1.32652f
C429 a_1198_518# a_1530_518# 0.307869f
C430 a_7718_4786# level_shifter_0.outb_h 0.183562f
C431 avss a_3854_518# 0.184675f
C432 avss a_2924_4788# 0.868706f
C433 avss ena 1.15253f
C434 avdd a_11138_9768# 0.071412f
C435 a_5862_4788# a_5704_4788# 0.036877f
C436 a_1842_9768# a_1510_9768# 0.307869f
C437 a_1012_7168# a_680_7168# 0.307869f
C438 avss a_7008_3118# 0.54635f
C439 avss a_9166_518# 0.184675f
C440 avss a_7154_9768# 0.142763f
C441 a_4036_4788# level_shifter_0.out_h 0.001601f
C442 avss a_846_9768# 0.142763f
C443 a_8482_9768# a_8150_9768# 0.307869f
C444 a_8336_3118# a_8004_3118# 0.307869f
C445 avdd a_11324_3118# 0.009316f
C446 avss a_4498_9768# 0.142763f
C447 level_shifter_0.outb_h a_6260_4788# 0.018927f
C448 avdd dout 0.101166f
C449 a_11636_7168# dvdd 1.06568f
C450 a_7672_3118# a_8004_3118# 0.307869f
C451 avss a_5470_5653# 0.001818f
C452 a_4830_9768# a_5162_9768# 0.307869f
C453 a_4166_9768# a_4498_9768# 0.307869f
C454 a_11636_7168# ena 0.098481f
C455 avdd a_9810_9768# 0.071412f
C456 a_1676_7168# a_2008_7168# 0.307869f
C457 avss a_11138_9768# 0.142763f
C458 avdd a_3336_7168# 0.548273f
C459 avdd a_1676_7168# 0.051033f
C460 avdd a_534_518# 0.031738f
C461 a_8980_7168# a_9312_7168# 0.307869f
C462 a_8714_4659# level_shifter_0.out_h 0.326647f
C463 a_3170_9768# a_2838_9768# 0.307869f
C464 a_4996_7168# a_5328_7168# 0.307869f
C465 avdd a_6490_9768# 0.071412f
C466 a_3688_3118# a_3356_3118# 0.307869f
C467 avdd a_4854_5653# 0.680997f
C468 avss a_11324_3118# 0.20921f
C469 a_5660_7168# a_5328_7168# 0.307869f
C470 avss dout 0.003814f
C471 a_4518_518# a_4850_518# 0.307869f
C472 a_7652_7168# a_7984_7168# 0.307869f
C473 level_shifter_0.inb_l a_9644_7168# 2.07e-20
C474 a_3006_5653# a_2924_4788# 4.31e-20
C475 a_6086_5653# a_6702_5653# 0.00665f
C476 a_1364_3118# a_1696_3118# 0.307869f
C477 avdd a_2838_9768# 0.071412f
C478 avss a_9810_9768# 0.142763f
C479 a_7718_4786# a_8714_4659# 0.007088f
C480 avdd a_6822_9768# 0.071412f
C481 avss a_3336_7168# 0.209517f
C482 avss a_1676_7168# 0.228829f
C483 avdd a_6842_518# 0.012005f
C484 avss a_534_518# 0.348434f
C485 a_11636_7168# a_11324_3118# 0.325625f
C486 a_8170_518# a_8502_518# 0.307869f
C487 a_11636_7168# dout 0.059654f
C488 avdd a_3622_5653# 0.790633f
C489 a_8668_3118# level_shifter_0.out_h 3.05e-19
C490 avss a_6490_9768# 0.142763f
C491 avdd a_680_7168# 0.055351f
C492 avss a_4854_5653# 0.002325f
C493 a_5862_4788# a_6086_5653# 0.015874f
C494 a_6344_3118# avss 0.739782f
C495 a_1842_9768# a_2174_9768# 0.307869f
C496 avdd a_9478_9768# 0.071412f
C497 avss a_7340_3118# 0.348693f
C498 a_5862_4788# level_shifter_0.out_h 0.164806f
C499 a_6324_7168# a_5992_7168# 0.307869f
C500 avss a_2838_9768# 0.142763f
C501 avdd a_10660_3118# 0.009316f
C502 a_5182_518# a_4850_518# 0.307869f
C503 avdd a_8482_9768# 0.071412f
C504 avdd a_4996_7168# 0.075453f
C505 level_shifter_0.inb_l level_shifter_0.outb_h 0.228327f
C506 a_9146_9768# a_9478_9768# 0.307869f
C507 avdd a_514_7168# 0.825392f
C508 avdd a_5660_7168# 0.548273f
C509 avss a_6822_9768# 0.142763f
C510 a_5162_9768# a_5494_9768# 0.307869f
C511 a_10308_7168# a_9976_7168# 0.307869f
C512 avss a_3688_3118# 0.353257f
C513 dvdd ena 1.57004f
C514 a_5826_9768# a_5494_9768# 0.307869f
C515 avss a_6842_518# 0.184675f
C516 avdd a_3668_7168# 0.548273f
C517 avss a_5704_4788# 0.86884f
C518 a_5862_4788# a_7718_4786# 4.61e-21
C519 a_10826_518# avdd 0.012005f
C520 avss a_5016_3118# 0.39682f
C521 a_7818_9768# a_8150_9768# 0.307869f
C522 avss a_680_7168# 0.238959f
C523 a_4684_3118# a_5016_3118# 0.307869f
C524 avdd a_7984_7168# 0.047956f
C525 avdd a_11890_5939# 6.58e-20
C526 avss a_9478_9768# 0.142763f
C527 avdd a_11304_7168# 0.516263f
C528 avdd a_4830_9768# 0.071412f
C529 a_5862_4788# a_6260_4788# 0.175672f
C530 avss a_8482_9768# 0.142763f
C531 avss a_10660_3118# 0.20921f
C532 avss a_4996_7168# 0.209517f
C533 avss a_514_7168# 2.39958f
C534 avss a_5660_7168# 0.209517f
C535 a_10826_518# a_11158_518# 0.307869f
C536 avdd a_10308_7168# 0.609955f
C537 avdd a_9332_3118# 0.032475f
C538 avdd a_9482_5327# 0.528099f
C539 a_8336_3118# a_8668_3118# 0.307869f
C540 a_7174_518# a_6842_518# 0.307869f
C541 a_866_518# a_1198_518# 0.307869f
C542 avss a_3668_7168# 0.209517f
C543 a_10826_518# avss 0.184675f
C544 dout dvss 1.18563f
C545 ena dvss 1.822f
C546 dvdd dvss 6.22115f
C547 avss dvss 6.815358f
C548 avdd dvss 0.392133p
C549 a_11490_518# dvss 0.297186f
C550 a_11324_3118# dvss 0.241933f
C551 a_11158_518# dvss 0.261223f
C552 a_10992_3118# dvss 0.241933f
C553 a_10826_518# dvss 0.261223f
C554 a_10660_3118# dvss 0.241933f
C555 a_10494_518# dvss 0.261223f
C556 a_10328_3118# dvss 0.254752f
C557 a_10162_518# dvss 0.261223f
C558 a_9996_3118# dvss 0.255929f
C559 a_9830_518# dvss 0.261223f
C560 a_9664_3118# dvss 0.241933f
C561 a_9498_518# dvss 0.261223f
C562 a_9332_3118# dvss 0.241933f
C563 a_9166_518# dvss 0.261223f
C564 a_9000_3118# dvss 0.241933f
C565 a_8834_518# dvss 0.261223f
C566 a_8668_3118# dvss 0.241933f
C567 a_8502_518# dvss 0.261223f
C568 a_8336_3118# dvss 0.241933f
C569 a_8170_518# dvss 0.261223f
C570 a_8004_3118# dvss 0.241933f
C571 a_7838_518# dvss 0.261223f
C572 a_7672_3118# dvss 0.241933f
C573 a_7506_518# dvss 0.261223f
C574 a_7340_3118# dvss 0.241933f
C575 a_7174_518# dvss 0.261223f
C576 a_7008_3118# dvss 0.241933f
C577 a_6842_518# dvss 0.261223f
C578 a_6676_3118# dvss 0.241933f
C579 a_6510_518# dvss 0.261223f
C580 a_6344_3118# dvss 0.241933f
C581 a_6178_518# dvss 0.261223f
C582 a_6012_3118# dvss 0.241933f
C583 a_5846_518# dvss 0.261223f
C584 a_5680_3118# dvss 0.241933f
C585 a_5514_518# dvss 0.261223f
C586 a_5348_3118# dvss 0.241933f
C587 a_5182_518# dvss 0.261223f
C588 a_5016_3118# dvss 0.241933f
C589 a_4850_518# dvss 0.261223f
C590 a_4684_3118# dvss 0.241933f
C591 a_4518_518# dvss 0.261223f
C592 a_4352_3118# dvss 0.241933f
C593 a_4186_518# dvss 0.261223f
C594 a_4020_3118# dvss 0.241933f
C595 a_3854_518# dvss 0.261223f
C596 a_3688_3118# dvss 0.241933f
C597 a_3522_518# dvss 0.261223f
C598 a_3356_3118# dvss 0.241933f
C599 a_3190_518# dvss 0.261223f
C600 a_3024_3118# dvss 0.241933f
C601 a_2858_518# dvss 0.261223f
C602 a_2692_3118# dvss 0.241933f
C603 a_2526_518# dvss 0.261223f
C604 a_2360_3118# dvss 0.241933f
C605 a_2194_518# dvss 0.261223f
C606 a_2028_3118# dvss 0.241933f
C607 a_1862_518# dvss 0.261223f
C608 a_1696_3118# dvss 0.241933f
C609 a_1530_518# dvss 0.261223f
C610 a_1364_3118# dvss 0.241933f
C611 a_1198_518# dvss 0.261223f
C612 a_1032_3118# dvss 0.24439f
C613 a_866_518# dvss 0.261223f
C614 a_700_3118# dvss 0.249183f
C615 a_534_518# dvss 0.296272f
C616 a_11890_5939# dvss 0.633389f
C617 a_7560_4786# dvss 0.011095f
C618 a_6260_4788# dvss 0.00951f
C619 a_5704_4788# dvss 0.00951f
C620 a_5148_4788# dvss 0.00951f
C621 a_4592_4788# dvss 0.00951f
C622 a_4036_4788# dvss 0.00951f
C623 a_3480_4788# dvss 0.00951f
C624 a_2924_4788# dvss 0.011998f
C625 a_2526_4188# dvss 0.00951f
C626 a_9482_5327# dvss 0.008785f
C627 a_8714_4659# dvss 0.008559f
C628 level_shifter_0.outb_h dvss 5.057272f
C629 level_shifter_0.inb_l dvss 0.970466f
C630 a_7718_4786# dvss 0.857037f
C631 a_5862_4788# dvss 0.146786f
C632 level_shifter_0.out_h dvss 5.442275f
C633 a_6702_5653# dvss 0.00886f
C634 a_6086_5653# dvss 0.00886f
C635 a_5470_5653# dvss 0.00886f
C636 a_4854_5653# dvss 0.00886f
C637 a_4238_5653# dvss 0.00886f
C638 a_3622_5653# dvss 0.00886f
C639 a_3006_5653# dvss 0.00886f
C640 a_11636_7168# dvss 2.90914f
C641 a_11470_9768# dvss 0.296245f
C642 a_11304_7168# dvss 0.241107f
C643 a_11138_9768# dvss 0.261295f
C644 a_10972_7168# dvss 0.240839f
C645 a_10806_9768# dvss 0.261295f
C646 a_10640_7168# dvss 0.240839f
C647 a_10474_9768# dvss 0.261295f
C648 a_10308_7168# dvss 0.240839f
C649 a_10142_9768# dvss 0.261295f
C650 a_9976_7168# dvss 0.240839f
C651 a_9810_9768# dvss 0.261295f
C652 a_9644_7168# dvss 0.242958f
C653 a_9478_9768# dvss 0.261295f
C654 a_9312_7168# dvss 0.240839f
C655 a_9146_9768# dvss 0.261295f
C656 a_8980_7168# dvss 0.240839f
C657 a_8814_9768# dvss 0.261295f
C658 a_8648_7168# dvss 0.240839f
C659 a_8482_9768# dvss 0.261295f
C660 a_8316_7168# dvss 0.240839f
C661 a_8150_9768# dvss 0.261295f
C662 a_7984_7168# dvss 0.240839f
C663 a_7818_9768# dvss 0.261295f
C664 a_7652_7168# dvss 0.240839f
C665 a_7486_9768# dvss 0.261295f
C666 a_7320_7168# dvss 0.240839f
C667 a_7154_9768# dvss 0.261295f
C668 a_6988_7168# dvss 0.240839f
C669 a_6822_9768# dvss 0.261295f
C670 a_6656_7168# dvss 0.240839f
C671 a_6490_9768# dvss 0.261295f
C672 a_6324_7168# dvss 0.240839f
C673 a_6158_9768# dvss 0.261295f
C674 a_5992_7168# dvss 0.240839f
C675 a_5826_9768# dvss 0.261295f
C676 a_5660_7168# dvss 0.240839f
C677 a_5494_9768# dvss 0.261295f
C678 a_5328_7168# dvss 0.240839f
C679 a_5162_9768# dvss 0.261295f
C680 a_4996_7168# dvss 0.240839f
C681 a_4830_9768# dvss 0.261295f
C682 a_4664_7168# dvss 0.240839f
C683 a_4498_9768# dvss 0.261295f
C684 a_4332_7168# dvss 0.240839f
C685 a_4166_9768# dvss 0.261295f
C686 a_4000_7168# dvss 0.240839f
C687 a_3834_9768# dvss 0.261295f
C688 a_3668_7168# dvss 0.240839f
C689 a_3502_9768# dvss 0.261295f
C690 a_3336_7168# dvss 0.240839f
C691 a_3170_9768# dvss 0.261295f
C692 a_3004_7168# dvss 0.240839f
C693 a_2838_9768# dvss 0.261295f
C694 a_2672_7168# dvss 0.240839f
C695 a_2506_9768# dvss 0.261295f
C696 a_2340_7168# dvss 0.240839f
C697 a_2174_9768# dvss 0.261295f
C698 a_2008_7168# dvss 0.240839f
C699 a_1842_9768# dvss 0.261295f
C700 a_1676_7168# dvss 0.240839f
C701 a_1510_9768# dvss 0.261295f
C702 a_1344_7168# dvss 0.240839f
C703 a_1178_9768# dvss 0.261295f
C704 a_1012_7168# dvss 0.240839f
C705 a_846_9768# dvss 0.261295f
C706 a_680_7168# dvss 0.240839f
C707 a_514_7168# dvss 0.139902f
C708 a_514_9768# dvss 0.297362f
C709 a_2982_4700.n0 dvss 2.14348f
C710 a_2982_4700.t3 dvss 0.165851f
C711 a_2982_4700.t5 dvss 0.164149f
C712 a_2982_4700.t0 dvss 0.031056f
C713 a_2982_4700.t2 dvss 0.162716f
C714 a_2982_4700.t4 dvss 0.153424f
C715 a_2982_4700.n1 dvss 1.14864f
C716 a_2982_4700.t1 dvss 0.030681f
C717 a_5306_4788.t2 dvss 3.77108f
C718 a_5306_4788.t0 dvss 0.010462f
C719 a_5306_4788.t4 dvss 0.05214f
C720 a_5306_4788.t3 dvss 0.055981f
C721 a_5306_4788.t1 dvss 0.010341f
C722 a_1414_4786.n0 dvss 7.603701f
C723 a_1414_4786.t3 dvss 0.068384f
C724 a_1414_4786.t4 dvss 0.349517f
C725 a_1414_4786.t6 dvss 0.342485f
C726 a_1414_4786.t5 dvss 0.342485f
C727 a_1414_4786.t8 dvss 0.342485f
C728 a_1414_4786.t11 dvss 0.342485f
C729 a_1414_4786.t7 dvss 0.342485f
C730 a_1414_4786.t10 dvss 0.342485f
C731 a_1414_4786.t9 dvss 0.342485f
C732 a_1414_4786.t2 dvss 0.072347f
C733 a_1414_4786.t0 dvss 0.342485f
C734 a_1414_4786.t1 dvss 0.066175f
C735 a_4750_4788.t2 dvss 3.67145f
C736 a_4750_4788.t0 dvss 0.010376f
C737 a_4750_4788.t4 dvss 0.0521f
C738 a_4750_4788.t3 dvss 0.055743f
C739 a_4750_4788.t1 dvss 0.01033f
C740 a_3082_4788.t2 dvss 3.38258f
C741 a_3082_4788.t1 dvss 0.009367f
C742 a_3082_4788.t4 dvss 0.047852f
C743 a_3082_4788.t3 dvss 0.050719f
C744 a_3082_4788.t0 dvss 0.009487f
C745 level_shifter_0.out_h.n0 dvss 3.99803f
C746 level_shifter_0.out_h.t5 dvss 0.266754f
C747 level_shifter_0.out_h.t1 dvss 0.050519f
C748 level_shifter_0.out_h.t0 dvss 0.050397f
C749 level_shifter_0.out_h.t4 dvss 0.310921f
C750 level_shifter_0.out_h.t6 dvss 0.259169f
C751 level_shifter_0.out_h.t3 dvss 0.252779f
C752 level_shifter_0.out_h.t2 dvss 0.283777f
C753 level_shifter_0.outb_h.n0 dvss 2.27957f
C754 level_shifter_0.outb_h.t2 dvss 0.661159f
C755 level_shifter_0.outb_h.t0 dvss 0.050895f
C756 level_shifter_0.outb_h.t3 dvss 0.315276f
C757 level_shifter_0.outb_h.t1 dvss 0.051265f
C758 level_shifter_0.outb_h.t4 dvss 0.273065f
C759 avdd.n0 dvss 14.7255f
C760 avdd.n1 dvss 6.24147f
C761 avdd.n2 dvss 4.02618f
C762 avdd.n3 dvss 0.647206f
C763 avdd.t2 dvss 0.020288f
C764 avdd.n4 dvss 0.43971f
C765 avdd.t4 dvss 0.020288f
C766 avdd.n5 dvss 0.43971f
C767 avdd.t12 dvss 0.020288f
C768 avdd.n6 dvss 0.038735f
C769 avdd.n7 dvss 0.129043f
C770 avdd.n8 dvss 0.033495f
C771 avdd.n9 dvss 0.034251f
C772 avdd.n10 dvss 0.129043f
C773 avdd.n11 dvss 0.117923f
C774 avdd.n12 dvss 0.117853f
C775 avdd.n13 dvss 0.117853f
C776 avdd.n14 dvss 1.21523f
C777 avdd.n15 dvss 0.117923f
C778 avdd.n16 dvss 1.21523f
C779 avdd.n17 dvss 0.117853f
C780 avdd.n18 dvss 0.117853f
C781 avdd.n19 dvss 0.159126f
C782 avdd.n20 dvss 0.159126f
C783 avdd.n21 dvss 0.117853f
C784 avdd.n22 dvss 0.117853f
C785 avdd.n23 dvss 1.21523f
C786 avdd.n24 dvss 0.117923f
C787 avdd.n25 dvss 0.117923f
C788 avdd.n26 dvss 1.21523f
C789 avdd.n27 dvss 0.033495f
C790 avdd.n28 dvss 0.117853f
C791 avdd.n29 dvss 0.034251f
C792 avdd.n30 dvss 0.038735f
C793 avdd.n31 dvss 0.110532f
C794 avdd.n32 dvss 0.117853f
C795 avdd.n33 dvss 0.039485f
C796 avdd.n34 dvss 0.039485f
C797 avdd.n35 dvss 0.034251f
C798 avdd.n36 dvss 0.24939f
C799 avdd.n37 dvss 0.117853f
C800 avdd.n38 dvss 0.117853f
C801 avdd.n39 dvss 1.98116f
C802 avdd.n40 dvss 0.117923f
C803 avdd.n41 dvss 1.21523f
C804 avdd.n42 dvss 0.117923f
C805 avdd.n43 dvss 0.117853f
C806 avdd.n44 dvss 0.117853f
C807 avdd.n45 dvss 0.502178f
C808 avdd.n46 dvss 0.034251f
C809 avdd.n47 dvss 1.12168f
C810 avdd.n48 dvss 1.09164f
C811 avdd.n49 dvss 0.117853f
C812 avdd.n50 dvss 0.317977f
C813 avdd.n51 dvss 0.24939f
C814 avdd.n52 dvss 0.276361f
C815 avdd.n53 dvss 0.117923f
C816 avdd.n55 dvss 1.97886f
C817 avdd.t23 dvss 1.52448f
C818 avdd.n56 dvss 0.117923f
C819 avdd.n57 dvss 0.131398f
C820 avdd.n58 dvss 0.339916f
C821 avdd.n59 dvss 0.038735f
C822 avdd.n60 dvss 0.340877f
C823 avdd.n61 dvss 0.039485f
C824 avdd.n62 dvss 0.129043f
C825 avdd.n63 dvss 0.110532f
C826 avdd.n64 dvss 0.038735f
C827 avdd.n65 dvss 0.213195f
C828 avdd.n66 dvss 0.229131f
C829 avdd.n67 dvss 0.033495f
C830 avdd.n68 dvss 0.159126f
C831 avdd.n69 dvss 0.150622f
C832 avdd.n70 dvss 0.117923f
C833 avdd.t3 dvss 1.28459f
C834 avdd.n71 dvss 0.117923f
C835 avdd.n72 dvss 0.150622f
C836 avdd.n73 dvss 0.15958f
C837 avdd.n74 dvss 0.15958f
C838 avdd.n75 dvss 0.150622f
C839 avdd.n76 dvss 0.15958f
C840 avdd.n77 dvss 0.15958f
C841 avdd.n78 dvss 0.150622f
C842 avdd.n79 dvss 0.15958f
C843 avdd.n80 dvss 0.15958f
C844 avdd.n81 dvss 0.117923f
C845 avdd.n82 dvss 0.117923f
C846 avdd.t13 dvss 1.28459f
C847 avdd.n83 dvss 0.117923f
C848 avdd.n84 dvss 0.033495f
C849 avdd.n85 dvss 0.117853f
C850 avdd.n86 dvss 0.117853f
C851 avdd.t5 dvss 1.28459f
C852 avdd.n87 dvss 0.117923f
C853 avdd.n88 dvss 0.117923f
C854 avdd.n89 dvss 0.131547f
C855 avdd.n90 dvss 1.53626f
C856 avdd.n91 dvss 0.102891f
C857 avdd.n92 dvss 0.159126f
C858 avdd.n93 dvss 0.159126f
C859 avdd.t6 dvss 0.020288f
C860 avdd.n94 dvss 0.43971f
C861 avdd.n95 dvss 0.129043f
C862 avdd.n96 dvss 0.150622f
C863 avdd.n97 dvss 0.039485f
C864 avdd.n98 dvss 0.15958f
C865 avdd.n99 dvss 0.117923f
C866 avdd.n100 dvss 0.034251f
C867 avdd.n101 dvss 1.21523f
C868 avdd.n102 dvss 0.150622f
C869 avdd.n103 dvss 0.159126f
C870 avdd.n104 dvss 0.110532f
C871 avdd.n105 dvss 0.038735f
C872 avdd.t10 dvss 0.020288f
C873 avdd.n106 dvss 0.43971f
C874 avdd.n107 dvss 0.110532f
C875 avdd.n108 dvss 0.15958f
C876 avdd.n109 dvss 0.117923f
C877 avdd.n110 dvss 0.117853f
C878 avdd.n111 dvss 0.150622f
C879 avdd.n112 dvss 1.21523f
C880 avdd.n113 dvss 0.117923f
C881 avdd.n114 dvss 0.117853f
C882 avdd.n115 dvss 0.117853f
C883 avdd.n116 dvss 0.159126f
C884 avdd.n117 dvss 0.033495f
C885 avdd.n118 dvss 0.038735f
C886 avdd.n119 dvss 0.159126f
C887 avdd.n120 dvss 0.117853f
C888 avdd.n121 dvss 0.117853f
C889 avdd.n122 dvss 1.21523f
C890 avdd.n123 dvss 0.117923f
C891 avdd.n124 dvss 0.117923f
C892 avdd.n125 dvss 1.21523f
C893 avdd.n126 dvss 0.129043f
C894 avdd.n127 dvss 0.033495f
C895 avdd.n128 dvss 0.117853f
C896 avdd.n129 dvss 0.034251f
C897 avdd.n130 dvss 0.038735f
C898 avdd.n131 dvss 0.129043f
C899 avdd.t16 dvss 0.020288f
C900 avdd.n132 dvss 0.697801f
C901 avdd.n133 dvss 2.47812f
C902 avdd.t8 dvss 0.020288f
C903 avdd.n134 dvss 0.117853f
C904 avdd.n135 dvss 0.039485f
C905 avdd.n136 dvss 0.039485f
C906 avdd.n137 dvss 0.258369f
C907 avdd.n138 dvss 0.117853f
C908 avdd.n139 dvss 0.117853f
C909 avdd.n140 dvss 1.21523f
C910 avdd.n141 dvss 0.117923f
C911 avdd.n142 dvss 1.21523f
C912 avdd.n143 dvss 0.117923f
C913 avdd.n144 dvss 0.117853f
C914 avdd.n145 dvss 0.117853f
C915 avdd.n146 dvss 0.159126f
C916 avdd.n147 dvss 0.117483f
C917 avdd.n148 dvss 0.082067f
C918 avdd.n149 dvss 0.132841f
C919 avdd.n150 dvss 0.281809f
C920 avdd.n151 dvss 0.080719f
C921 avdd.n152 dvss 0.255802f
C922 avdd.n153 dvss 0.247546f
C923 avdd.n154 dvss 0.117923f
C924 avdd.t15 dvss 1.28459f
C925 avdd.n155 dvss 0.117923f
C926 avdd.n156 dvss 0.249297f
C927 avdd.n157 dvss 0.15958f
C928 avdd.n158 dvss 0.15958f
C929 avdd.n159 dvss 0.150622f
C930 avdd.n160 dvss 0.15958f
C931 avdd.n161 dvss 0.15958f
C932 avdd.n162 dvss 0.034251f
C933 avdd.n163 dvss 0.229131f
C934 avdd.n164 dvss 0.213195f
C935 avdd.n165 dvss 0.43971f
C936 avdd.n166 dvss 1.15036f
C937 avdd.t18 dvss 0.0203f
C938 avdd.n167 dvss 0.590731f
C939 avdd.n168 dvss 0.213195f
C940 avdd.n169 dvss 0.229131f
C941 avdd.n170 dvss 0.110532f
C942 avdd.n171 dvss 0.117923f
C943 avdd.t7 dvss 1.28459f
C944 avdd.n172 dvss 0.117923f
C945 avdd.n173 dvss 0.150622f
C946 avdd.n174 dvss 0.159126f
C947 avdd.n175 dvss 0.159126f
C948 avdd.n176 dvss 0.150622f
C949 avdd.n177 dvss 0.117923f
C950 avdd.t9 dvss 1.28459f
C951 avdd.n178 dvss 0.117923f
C952 avdd.n179 dvss 0.117853f
C953 avdd.n180 dvss 0.039485f
C954 avdd.n181 dvss 0.129043f
C955 avdd.n182 dvss 0.213195f
C956 avdd.n183 dvss 0.229131f
C957 avdd.n184 dvss 0.033495f
C958 avdd.n185 dvss 0.117853f
C959 avdd.n186 dvss 1.21523f
C960 avdd.n187 dvss 0.117853f
C961 avdd.n188 dvss 0.117923f
C962 avdd.n189 dvss 0.150622f
C963 avdd.n190 dvss 0.15958f
C964 avdd.n191 dvss 0.15958f
C965 avdd.n192 dvss 0.034251f
C966 avdd.n193 dvss 0.229131f
C967 avdd.n194 dvss 0.213195f
C968 avdd.n195 dvss 0.038735f
C969 avdd.n196 dvss 0.117853f
C970 avdd.n197 dvss 1.21523f
C971 avdd.n198 dvss 1.21523f
C972 avdd.n199 dvss 0.117853f
C973 avdd.n200 dvss 0.117923f
C974 avdd.n201 dvss 0.117853f
C975 avdd.n202 dvss 1.21523f
C976 avdd.n203 dvss 0.117853f
C977 avdd.n204 dvss 0.039485f
C978 avdd.n205 dvss 0.129043f
C979 avdd.t14 dvss 0.020288f
C980 avdd.n206 dvss 0.43971f
C981 avdd.n207 dvss 0.213195f
C982 avdd.n208 dvss 0.229131f
C983 avdd.n209 dvss 0.110532f
C984 avdd.n210 dvss 0.117923f
C985 avdd.t11 dvss 1.28459f
C986 avdd.n211 dvss 0.117923f
C987 avdd.n212 dvss 0.150622f
C988 avdd.n213 dvss 0.159126f
C989 avdd.n214 dvss 0.159126f
C990 avdd.n215 dvss 0.150622f
C991 avdd.n216 dvss 0.117923f
C992 avdd.t1 dvss 1.28459f
C993 avdd.n217 dvss 0.117923f
C994 avdd.n218 dvss 0.110532f
C995 avdd.n219 dvss 0.229131f
C996 avdd.n220 dvss 0.213195f
C997 avdd.n221 dvss 0.43971f
C998 avdd.n222 dvss 1.15036f
C999 avdd.n223 dvss 2.74093f
C1000 avdd.n224 dvss 5.46532f
C1001 avdd.n225 dvss 2.78737f
C1002 avdd.n226 dvss 6.01336f
C1003 avdd.n227 dvss 1.08997f
C1004 avdd.n228 dvss 3.15497f
C1005 avdd.n229 dvss 0.904845f
C1006 avdd.n230 dvss 13.5245f
C1007 avdd.n231 dvss 2.97694f
C1008 avdd.n232 dvss 1.63592f
C1009 avdd.n233 dvss 0.743661f
C1010 avdd.n234 dvss 0.117923f
C1011 avdd.n235 dvss 0.117923f
C1012 avdd.n236 dvss 0.30969f
C1013 avdd.n237 dvss 0.13157f
C1014 avdd.n238 dvss 0.98242f
C1015 avdd.n239 dvss 2.48826f
C1016 avdd.n240 dvss 3.15514f
C1017 avdd.n241 dvss 4.47652f
C1018 avdd.n242 dvss 3.202f
C1019 avdd.n243 dvss 3.70777f
C1020 avdd.n244 dvss 16.0032f
C1021 avdd.n245 dvss 13.5252f
C1022 avdd.n246 dvss 7.71493f
C1023 avdd.n247 dvss 1.80014f
C1024 avdd.n248 dvss 0.904682f
C1025 avdd.n249 dvss 1.50347f
C1026 avdd.n250 dvss 0.855737f
C1027 avdd.n251 dvss 0.737356f
C1028 avdd.n252 dvss 1.33731f
C1029 avdd.t20 dvss 0.020263f
C1030 avdd.n253 dvss 0.258583f
C1031 avdd.t22 dvss 0.020263f
C1032 avdd.n254 dvss 0.124128f
C1033 avdd.n255 dvss 0.236114f
C1034 avdd.n256 dvss 0.117853f
C1035 avdd.n257 dvss 0.117853f
C1036 avdd.n258 dvss 1.38607f
C1037 avdd.n259 dvss 0.117923f
C1038 avdd.n260 dvss 0.117923f
C1039 avdd.n261 dvss 1.40702f
C1040 avdd.n262 dvss 0.568074f
C1041 avdd.n263 dvss 0.179944f
C1042 avdd.n264 dvss 0.117923f
C1043 avdd.n265 dvss 0.215466f
C1044 avdd.n266 dvss 0.117853f
C1045 avdd.n267 dvss 0.123732f
C1046 avdd.n268 dvss 0.093275f
C1047 avdd.n269 dvss 0.117923f
C1048 avdd.t19 dvss 0.743661f
C1049 avdd.t21 dvss 0.743661f
C1050 avdd.n270 dvss 0.142964f
C1051 avdd.n271 dvss 0.243088f
C1052 avdd.n272 dvss 0.117853f
C1053 avdd.n273 dvss 0.743661f
C1054 avdd.n274 dvss 0.663359f
C1055 avdd.n275 dvss 0.117853f
C1056 avdd.n276 dvss 0.110532f
C1057 avdd.n277 dvss 0.117853f
C1058 avdd.n278 dvss 0.135256f
C1059 avdd.n279 dvss 0.28079f
C1060 avdd.n280 dvss 0.177629f
C1061 avdd.n281 dvss 0.117853f
C1062 avdd.n282 dvss 0.208845f
C1063 avdd.n283 dvss 0.308299f
C1064 avdd.n284 dvss 0.214712f
C1065 avdd.n285 dvss 0.117923f
C1066 avdd.t17 dvss 1.48184f
C1067 avdd.n286 dvss 0.117923f
C1068 avdd.n287 dvss 0.13474f
C1069 avdd.n288 dvss 0.158253f
C1070 avdd.n289 dvss -0.071355f
C1071 avdd.n290 dvss -2.12191f
C1072 avdd.n291 dvss 1.66562f
C1073 avdd.n292 dvss 0.160339f
C1074 avdd.n293 dvss 0.127531f
C1075 avdd.n294 dvss 0.117853f
C1076 avdd.n295 dvss 0.991547f
C1077 avdd.n296 dvss 3.96545f
C1078 avdd.n297 dvss 3.69809f
C1079 avdd.n298 dvss 7.71766f
C1080 avdd.n299 dvss 1.8008f
C1081 avdd.n300 dvss 0.633609f
C1082 avdd.n301 dvss 2.34564f
C1083 avdd.n302 dvss 7.20856f
C1084 avdd.n303 dvss 31.262098f
C1085 avdd.n304 dvss 36.207603f
C1086 avdd.n305 dvss 30.1327f
C1087 avdd.n306 dvss 18.317598f
C1088 a_2368_4788.n0 dvss 4.61781f
C1089 a_2368_4788.n1 dvss 1.89182f
C1090 a_2368_4788.t0 dvss 0.32443f
C1091 a_2368_4788.t7 dvss 0.32443f
C1092 a_2368_4788.t6 dvss 0.32443f
C1093 a_2368_4788.t8 dvss 0.32443f
C1094 a_2368_4788.t4 dvss 0.32443f
C1095 a_2368_4788.t5 dvss 0.32443f
C1096 a_2368_4788.t10 dvss 0.32443f
C1097 a_2368_4788.t9 dvss 0.331908f
C1098 a_2368_4788.t3 dvss 0.064406f
C1099 a_2368_4788.t2 dvss 0.061523f
C1100 a_2368_4788.t1 dvss 0.061523f
C1101 a_4194_4788.t4 dvss 3.57109f
C1102 a_4194_4788.t1 dvss 0.010379f
C1103 a_4194_4788.t3 dvss 0.052339f
C1104 a_4194_4788.t2 dvss 0.055811f
C1105 a_4194_4788.t0 dvss 0.010378f
C1106 a_3638_4788.t3 dvss 3.57257f
C1107 a_3638_4788.t0 dvss 0.010209f
C1108 a_3638_4788.t2 dvss 0.05184f
C1109 a_3638_4788.t4 dvss 0.055102f
C1110 a_3638_4788.t1 dvss 0.010278f
C1111 avss.n0 dvss 6.17475f
C1112 avss.n1 dvss 1.35168f
C1113 avss.n2 dvss 1.94176f
C1114 avss.n3 dvss 0.58426f
C1115 avss.n4 dvss 0.58426f
C1116 avss.t124 dvss 0.619705f
C1117 avss.n5 dvss 0.060862f
C1118 avss.n6 dvss 0.060862f
C1119 avss.n7 dvss 0.146424f
C1120 avss.n8 dvss 0.071574f
C1121 avss.t51 dvss 0.010452f
C1122 avss.n9 dvss 0.234041f
C1123 avss.n10 dvss 0.13808f
C1124 avss.n11 dvss 1.99881f
C1125 avss.n12 dvss 10.249599f
C1126 avss.t139 dvss 0.010342f
C1127 avss.n13 dvss 0.066335f
C1128 avss.n14 dvss 0.01734f
C1129 avss.n15 dvss 0.01734f
C1130 avss.n16 dvss 0.01738f
C1131 avss.n17 dvss 0.01734f
C1132 avss.n18 dvss 0.060862f
C1133 avss.t92 dvss 0.010344f
C1134 avss.n19 dvss 0.174915f
C1135 avss.n20 dvss 0.040456f
C1136 avss.n21 dvss 0.060994f
C1137 avss.n22 dvss 0.060994f
C1138 avss.t40 dvss 1.25712f
C1139 avss.n23 dvss 0.060862f
C1140 avss.t145 dvss 1.11547f
C1141 avss.n24 dvss 0.072933f
C1142 avss.n25 dvss 0.01738f
C1143 avss.n26 dvss 0.073499f
C1144 avss.t117 dvss 1.12137f
C1145 avss.n27 dvss 0.908901f
C1146 avss.t90 dvss 1.25028f
C1147 avss.n28 dvss 0.58426f
C1148 avss.n29 dvss 0.58426f
C1149 avss.n30 dvss 1.94031f
C1150 avss.n31 dvss 1.85919f
C1151 avss.n32 dvss 0.36127f
C1152 avss.t151 dvss 0.010318f
C1153 avss.n33 dvss 0.201702f
C1154 avss.n34 dvss 0.306529f
C1155 avss.n35 dvss 0.398641f
C1156 avss.n36 dvss 1.9049f
C1157 avss.t105 dvss 1.35108f
C1158 avss.t53 dvss 1.3351f
C1159 avss.t31 dvss 1.3351f
C1160 avss.t99 dvss 1.3351f
C1161 avss.t82 dvss 1.3351f
C1162 avss.t14 dvss 1.3351f
C1163 avss.t56 dvss 1.3351f
C1164 avss.t109 dvss 1.3351f
C1165 avss.t122 dvss 1.3351f
C1166 avss.t157 dvss 1.3351f
C1167 avss.t158 dvss 1.3351f
C1168 avss.t144 dvss 1.33699f
C1169 avss.t116 dvss 1.43767f
C1170 avss.t29 dvss 1.43592f
C1171 avss.t81 dvss 1.43592f
C1172 avss.t1 dvss 1.43592f
C1173 avss.t161 dvss 1.31049f
C1174 avss.t39 dvss 1.43631f
C1175 avss.t154 dvss 1.43631f
C1176 avss.t30 dvss 1.43631f
C1177 avss.t123 dvss 1.43631f
C1178 avss.t15 dvss 1.43631f
C1179 avss.t46 dvss 1.43631f
C1180 avss.t43 dvss 1.43631f
C1181 avss.t44 dvss 1.43631f
C1182 avss.t106 dvss 1.43631f
C1183 avss.t121 dvss 1.43631f
C1184 avss.t164 dvss 1.43631f
C1185 avss.t28 dvss 1.43631f
C1186 avss.t0 dvss 1.43631f
C1187 avss.t12 dvss 1.43631f
C1188 avss.t49 dvss 1.43631f
C1189 avss.t136 dvss 1.43631f
C1190 avss.t118 dvss 1.43631f
C1191 avss.t163 dvss 1.43631f
C1192 avss.t48 dvss 1.43631f
C1193 avss.t11 dvss 1.43631f
C1194 avss.t64 dvss 1.43631f
C1195 avss.t147 dvss 1.43631f
C1196 avss.t159 dvss 1.43631f
C1197 avss.t38 dvss 1.43631f
C1198 avss.t114 dvss 1.43631f
C1199 avss.t25 dvss 1.43631f
C1200 avss.t126 dvss 1.43631f
C1201 avss.t143 dvss 1.07723f
C1202 avss.n37 dvss 0.718153f
C1203 avss.t94 dvss 1.07723f
C1204 avss.t111 dvss 1.43631f
C1205 avss.t3 dvss 1.43631f
C1206 avss.t85 dvss 1.43631f
C1207 avss.t42 dvss 1.43631f
C1208 avss.t9 dvss 1.43632f
C1209 avss.t165 dvss 1.43593f
C1210 avss.t19 dvss 1.43592f
C1211 avss.t91 dvss 1.43592f
C1212 avss.t83 dvss 1.43592f
C1213 avss.t62 dvss 1.43592f
C1214 avss.t152 dvss 1.43592f
C1215 avss.t76 dvss 1.43592f
C1216 avss.t96 dvss 1.43592f
C1217 avss.t13 dvss 1.43592f
C1218 avss.t104 dvss 1.43592f
C1219 avss.t119 dvss 0.843384f
C1220 avss.n38 dvss 0.968429f
C1221 avss.n39 dvss 0.060862f
C1222 avss.n40 dvss 0.060862f
C1223 avss.n41 dvss 0.059005f
C1224 avss.n42 dvss 0.090237f
C1225 avss.n43 dvss 0.153956f
C1226 avss.n44 dvss 0.544628f
C1227 avss.n45 dvss 0.060994f
C1228 avss.t59 dvss 0.010352f
C1229 avss.n46 dvss 0.904763f
C1230 avss.n47 dvss 0.104788f
C1231 avss.t150 dvss 0.313974f
C1232 avss.t103 dvss 1.64296f
C1233 avss.n48 dvss 0.061012f
C1234 avss.t112 dvss 1.02694f
C1235 avss.n49 dvss 0.060862f
C1236 avss.n50 dvss 0.060862f
C1237 avss.n51 dvss 0.133072f
C1238 avss.n52 dvss 0.0173f
C1239 avss.n53 dvss 0.531478f
C1240 avss.n54 dvss 0.060994f
C1241 avss.t155 dvss 1.2099f
C1242 avss.n55 dvss 0.060862f
C1243 avss.n56 dvss 0.060994f
C1244 avss.t20 dvss 1.19219f
C1245 avss.n57 dvss 0.060862f
C1246 avss.n58 dvss 0.060862f
C1247 avss.n59 dvss 0.01734f
C1248 avss.n60 dvss 0.776783f
C1249 avss.n61 dvss 0.076242f
C1250 avss.n62 dvss 0.060862f
C1251 avss.n63 dvss 0.057388f
C1252 avss.t160 dvss 0.011239f
C1253 avss.n64 dvss 0.407008f
C1254 avss.n65 dvss 0.666495f
C1255 avss.t73 dvss 0.010342f
C1256 avss.n66 dvss 0.066335f
C1257 avss.n67 dvss 0.01734f
C1258 avss.n68 dvss 0.01734f
C1259 avss.n69 dvss 0.01734f
C1260 avss.n70 dvss 0.01734f
C1261 avss.n71 dvss 0.060862f
C1262 avss.n72 dvss 0.040955f
C1263 avss.n73 dvss 0.060994f
C1264 avss.n74 dvss 0.060994f
C1265 avss.t87 dvss 1.25712f
C1266 avss.n75 dvss 0.060862f
C1267 avss.t142 dvss 1.2099f
C1268 avss.n76 dvss 0.072589f
C1269 avss.n77 dvss 0.01734f
C1270 avss.n78 dvss 0.01734f
C1271 avss.n79 dvss 0.072589f
C1272 avss.n80 dvss 0.060994f
C1273 avss.n81 dvss 0.060994f
C1274 avss.t132 dvss 1.09186f
C1275 avss.n82 dvss 0.060862f
C1276 avss.n83 dvss 0.060862f
C1277 avss.t153 dvss 1.25712f
C1278 avss.n84 dvss 0.082768f
C1279 avss.n85 dvss 0.01734f
C1280 avss.n86 dvss 0.057388f
C1281 avss.t72 dvss 0.010342f
C1282 avss.n87 dvss 0.174138f
C1283 avss.n88 dvss 0.285735f
C1284 avss.n89 dvss 0.308497f
C1285 avss.t35 dvss 0.010342f
C1286 avss.n90 dvss 0.066335f
C1287 avss.n91 dvss 0.01734f
C1288 avss.n92 dvss 0.01734f
C1289 avss.n93 dvss 0.01734f
C1290 avss.n94 dvss 0.01734f
C1291 avss.n95 dvss 0.060862f
C1292 avss.n96 dvss 0.040955f
C1293 avss.n97 dvss 0.060994f
C1294 avss.n98 dvss 0.060994f
C1295 avss.t63 dvss 1.25712f
C1296 avss.n99 dvss 0.060862f
C1297 avss.t134 dvss 1.16269f
C1298 avss.n100 dvss 0.072589f
C1299 avss.n101 dvss 0.01734f
C1300 avss.n102 dvss 0.01734f
C1301 avss.n103 dvss 0.072589f
C1302 avss.n104 dvss 0.060994f
C1303 avss.n105 dvss 0.060994f
C1304 avss.t146 dvss 1.13908f
C1305 avss.n106 dvss 0.060862f
C1306 avss.n107 dvss 0.060862f
C1307 avss.t7 dvss 1.25712f
C1308 avss.n108 dvss 0.082768f
C1309 avss.n109 dvss 0.01734f
C1310 avss.n110 dvss 0.01734f
C1311 avss.n111 dvss 0.01734f
C1312 avss.n112 dvss 0.01734f
C1313 avss.n113 dvss 0.057388f
C1314 avss.t37 dvss 1.07416f
C1315 avss.n114 dvss 0.060994f
C1316 avss.t47 dvss 1.09776f
C1317 avss.n115 dvss 0.885293f
C1318 avss.n116 dvss 0.861685f
C1319 avss.n117 dvss 0.060994f
C1320 avss.n118 dvss 0.01734f
C1321 avss.n119 dvss 0.072589f
C1322 avss.n120 dvss 0.060994f
C1323 avss.n121 dvss 0.060994f
C1324 avss.t41 dvss 1.25712f
C1325 avss.n122 dvss 0.060862f
C1326 avss.t125 dvss 1.25712f
C1327 avss.n123 dvss 0.060862f
C1328 avss.n124 dvss 0.01734f
C1329 avss.n125 dvss 0.057388f
C1330 avss.t66 dvss 1.02694f
C1331 avss.n126 dvss 0.060994f
C1332 avss.t21 dvss 1.14498f
C1333 avss.n127 dvss 0.932509f
C1334 avss.n128 dvss 0.81447f
C1335 avss.n129 dvss 0.060994f
C1336 avss.n130 dvss 0.01734f
C1337 avss.n131 dvss 0.072589f
C1338 avss.n132 dvss 0.060994f
C1339 avss.n133 dvss 0.060994f
C1340 avss.t23 dvss 1.25712f
C1341 avss.n134 dvss 0.060862f
C1342 avss.t162 dvss 1.25712f
C1343 avss.n135 dvss 0.060862f
C1344 avss.n136 dvss 0.060994f
C1345 avss.n137 dvss 0.060994f
C1346 avss.n138 dvss 0.979724f
C1347 avss.t129 dvss 0.767254f
C1348 avss.n139 dvss 0.979724f
C1349 avss.n140 dvss 0.060994f
C1350 avss.n141 dvss 0.01734f
C1351 avss.n142 dvss 0.082768f
C1352 avss.n143 dvss 0.01734f
C1353 avss.t135 dvss 1.25712f
C1354 avss.t98 dvss 1.04465f
C1355 avss.t69 dvss 0.979724f
C1356 avss.n144 dvss 0.060862f
C1357 avss.n145 dvss 0.122263f
C1358 avss.n146 dvss 0.130265f
C1359 avss.n147 dvss 0.211201f
C1360 avss.n148 dvss 0.211282f
C1361 avss.n149 dvss 0.07941f
C1362 avss.n150 dvss 0.072589f
C1363 avss.n151 dvss 0.01734f
C1364 avss.n152 dvss 0.060994f
C1365 avss.n153 dvss 0.979724f
C1366 avss.t93 dvss 0.619705f
C1367 avss.n154 dvss 0.637411f
C1368 avss.n155 dvss 0.489862f
C1369 avss.n156 dvss 0.060994f
C1370 avss.n157 dvss 0.01734f
C1371 avss.n158 dvss 0.072589f
C1372 avss.n159 dvss 0.072589f
C1373 avss.n160 dvss 0.072589f
C1374 avss.n161 dvss 0.07941f
C1375 avss.n162 dvss 0.060862f
C1376 avss.t16 dvss 0.979724f
C1377 avss.n163 dvss 0.060862f
C1378 avss.n164 dvss 0.07941f
C1379 avss.n165 dvss 0.072589f
C1380 avss.n166 dvss 0.072589f
C1381 avss.n167 dvss 0.07941f
C1382 avss.n168 dvss 0.072589f
C1383 avss.n169 dvss 0.072589f
C1384 avss.n170 dvss 0.07326f
C1385 avss.n171 dvss 2.64461f
C1386 avss.n172 dvss 0.792859f
C1387 avss.n173 dvss 0.039035f
C1388 avss.n174 dvss 0.01734f
C1389 avss.n175 dvss 0.060994f
C1390 avss.n176 dvss 0.979724f
C1391 avss.t148 dvss 0.767254f
C1392 avss.n177 dvss 0.979724f
C1393 avss.n178 dvss 0.060994f
C1394 avss.n179 dvss 0.060994f
C1395 avss.n180 dvss 0.979724f
C1396 avss.t101 dvss 0.767254f
C1397 avss.n181 dvss 0.979724f
C1398 avss.n182 dvss 0.060994f
C1399 avss.n183 dvss 0.01734f
C1400 avss.n184 dvss 0.082768f
C1401 avss.n185 dvss 0.01734f
C1402 avss.n186 dvss 0.072589f
C1403 avss.n187 dvss 0.072589f
C1404 avss.n188 dvss 0.07941f
C1405 avss.n189 dvss 0.060862f
C1406 avss.t34 dvss 0.979724f
C1407 avss.n190 dvss 0.060862f
C1408 avss.n191 dvss 0.07941f
C1409 avss.n192 dvss 0.072589f
C1410 avss.n193 dvss 0.072589f
C1411 avss.n194 dvss 0.07941f
C1412 avss.n195 dvss 0.072589f
C1413 avss.n196 dvss 0.072589f
C1414 avss.n197 dvss 0.07941f
C1415 avss.n198 dvss 0.072589f
C1416 avss.n199 dvss 0.072589f
C1417 avss.n200 dvss 0.060862f
C1418 avss.n201 dvss 0.057118f
C1419 avss.n202 dvss 0.060994f
C1420 avss.n203 dvss 0.062984f
C1421 avss.n204 dvss 0.296871f
C1422 avss.n205 dvss 0.072589f
C1423 avss.n206 dvss 0.072589f
C1424 avss.n207 dvss 0.07941f
C1425 avss.n208 dvss 0.060862f
C1426 avss.n209 dvss 0.060994f
C1427 avss.n210 dvss 0.979724f
C1428 avss.t27 dvss 0.767254f
C1429 avss.t107 dvss 1.25712f
C1430 avss.n211 dvss 0.072589f
C1431 avss.n212 dvss 0.072573f
C1432 avss.n213 dvss 0.07941f
C1433 avss.n214 dvss 0.060862f
C1434 avss.n215 dvss 0.060994f
C1435 avss.n216 dvss 0.060994f
C1436 avss.n217 dvss 0.060994f
C1437 avss.n218 dvss 0.979724f
C1438 avss.t102 dvss 0.767254f
C1439 avss.n219 dvss 0.979724f
C1440 avss.t55 dvss 1.25712f
C1441 avss.t138 dvss 0.979724f
C1442 avss.n220 dvss 0.060862f
C1443 avss.n221 dvss 0.060994f
C1444 avss.n222 dvss 0.979724f
C1445 avss.n223 dvss 0.060994f
C1446 avss.n224 dvss 0.01734f
C1447 avss.n225 dvss 0.082768f
C1448 avss.n226 dvss 0.057388f
C1449 avss.t74 dvss 0.010342f
C1450 avss.n227 dvss 0.174138f
C1451 avss.n228 dvss 1.14995f
C1452 avss.n229 dvss 0.640978f
C1453 avss.n230 dvss 1.4189f
C1454 avss.t141 dvss 0.010342f
C1455 avss.n231 dvss 0.174138f
C1456 avss.n232 dvss 0.040955f
C1457 avss.n233 dvss 0.066335f
C1458 avss.n234 dvss 0.060862f
C1459 avss.t140 dvss 0.979724f
C1460 avss.n235 dvss 0.060862f
C1461 avss.n236 dvss 0.07941f
C1462 avss.n237 dvss 0.072589f
C1463 avss.n238 dvss 0.072589f
C1464 avss.n239 dvss 0.07941f
C1465 avss.n240 dvss 0.060862f
C1466 avss.t52 dvss 0.979724f
C1467 avss.n241 dvss 0.060862f
C1468 avss.n242 dvss 0.066335f
C1469 avss.n243 dvss 0.082768f
C1470 avss.n244 dvss 0.057388f
C1471 avss.n245 dvss 0.040955f
C1472 avss.n246 dvss 0.174138f
C1473 avss.n247 dvss 0.371066f
C1474 avss.n248 dvss 0.393726f
C1475 avss.t137 dvss 0.010342f
C1476 avss.n249 dvss 0.174138f
C1477 avss.n250 dvss 0.040955f
C1478 avss.n251 dvss 0.066335f
C1479 avss.n252 dvss 0.060862f
C1480 avss.t5 dvss 0.979724f
C1481 avss.n253 dvss 0.060862f
C1482 avss.n254 dvss 0.07941f
C1483 avss.n255 dvss 0.072589f
C1484 avss.n256 dvss 0.072589f
C1485 avss.n257 dvss 0.07941f
C1486 avss.n258 dvss 0.060862f
C1487 avss.t71 dvss 0.979724f
C1488 avss.n259 dvss 0.060862f
C1489 avss.n260 dvss 0.066335f
C1490 avss.n261 dvss 0.082768f
C1491 avss.n262 dvss 0.057388f
C1492 avss.n263 dvss 0.040955f
C1493 avss.n264 dvss 0.174138f
C1494 avss.n265 dvss 1.53575f
C1495 avss.n266 dvss 1.22337f
C1496 avss.n267 dvss 0.588805f
C1497 avss.n268 dvss 1.35874f
C1498 avss.t61 dvss 1.70171f
C1499 avss.t79 dvss 1.48535f
C1500 avss.t113 dvss 1.48535f
C1501 avss.t65 dvss 1.48535f
C1502 avss.t108 dvss 1.48535f
C1503 avss.t128 dvss 1.48535f
C1504 avss.t133 dvss 1.48535f
C1505 avss.t8 dvss 1.47754f
C1506 avss.t88 dvss 1.32856f
C1507 avss.t60 dvss 1.33355f
C1508 avss.t78 dvss 1.33355f
C1509 avss.t100 dvss 1.33355f
C1510 avss.t115 dvss 1.33355f
C1511 avss.t36 dvss 1.33355f
C1512 avss.t77 dvss 1.33355f
C1513 avss.t67 dvss 1.33355f
C1514 avss.t84 dvss 1.33355f
C1515 avss.t166 dvss 1.33355f
C1516 avss.t120 dvss 1.33355f
C1517 avss.t18 dvss 1.33933f
C1518 avss.n269 dvss 1.75287f
C1519 avss.n270 dvss 1.07463f
C1520 avss.n271 dvss 1.32864f
C1521 avss.n272 dvss 13.756599f
C1522 avss.n273 dvss 1.9833f
C1523 avss.t149 dvss 2.98637f
C1524 avss.n274 dvss 1.57997f
C1525 avss.t86 dvss 2.16856f
C1526 avss.n275 dvss 1.91931f
C1527 avss.t6 dvss 1.59974f
C1528 avss.n276 dvss 1.91916f
C1529 avss.t89 dvss 1.59974f
C1530 avss.t75 dvss 1.89088f
C1531 avss.n277 dvss 1.97303f
C1532 avss.n278 dvss 1.57954f
C1533 avss.n279 dvss 0.346192f
C1534 avss.n280 dvss 8.215039f
C1535 avss.n281 dvss 15.4977f
C1536 avss.n282 dvss 2.39644f
C1537 avss.t70 dvss 0.010342f
C1538 avss.n283 dvss 0.174138f
C1539 avss.n284 dvss 0.040955f
C1540 avss.n285 dvss 0.063067f
C1541 avss.n286 dvss 0.089331f
C1542 avss.n287 dvss 0.284185f
C1543 avss.n288 dvss 0.060994f
C1544 avss.n289 dvss 0.979724f
C1545 avss.t10 dvss 1.74698f
C1546 avss.t26 dvss 1.95945f
C1547 avss.t130 dvss 1.95945f
C1548 avss.t95 dvss 1.95945f
C1549 avss.t24 dvss 1.45188f
C1550 avss.n290 dvss 0.060994f
C1551 avss.n291 dvss 0.979724f
C1552 avss.t80 dvss 1.25712f
C1553 avss.t57 dvss 0.979724f
C1554 avss.n292 dvss 0.060862f
C1555 avss.n293 dvss 0.081601f
C1556 avss.n294 dvss 0.098331f
C1557 avss.n295 dvss 0.14206f
C1558 avss.n296 dvss 0.134005f
C1559 avss.n297 dvss 0.060994f
C1560 avss.n298 dvss 0.979724f
C1561 avss.t17 dvss 1.91223f
C1562 avss.t33 dvss 1.25121f
C1563 avss.n299 dvss 1.63635f
C1564 avss.n300 dvss 1.49568f
C1565 avss.n301 dvss 0.060994f
C1566 avss.n302 dvss 0.155039f
C1567 avss.n303 dvss 0.105179f
C1568 avss.n304 dvss 0.040092f
C1569 avss.n305 dvss 0.074707f
C1570 avss.n306 dvss 0.134148f
C1571 avss.n307 dvss 0.041649f
C1572 avss.n308 dvss 0.060862f
C1573 avss.t58 dvss 0.558778f
C1574 avss.n310 dvss 0.060862f
C1575 avss.n311 dvss 0.090792f
C1576 avss.n312 dvss 0.142421f
C1577 avss.n313 dvss 0.067616f
C1578 avss.n314 dvss 0.060994f
C1579 avss.n315 dvss 0.250473f
C1580 avss.n316 dvss 0.093212f
C1581 avss.n317 dvss 2.81827f
C1582 avss.n318 dvss 0.101659f
C1583 avss.n319 dvss 0.975596f
C1584 avss.n320 dvss 2.48839f
C1585 avss.n321 dvss 5.40126f
C1586 avss.n322 dvss 1.82062f
C1587 avss.t97 dvss 1.44742f
C1588 avss.t156 dvss 1.43631f
C1589 avss.t32 dvss 1.43631f
C1590 avss.t54 dvss 1.43631f
C1591 avss.t22 dvss 0.904181f
C1592 avss.n323 dvss 3.6879f
C1593 avss.n324 dvss 3.7429f
C1594 avss.t50 dvss 0.843979f
C1595 avss.t4 dvss 1.18629f
C1596 avss.t131 dvss 1.05055f
C1597 avss.n325 dvss 0.838078f
C1598 avss.n326 dvss 0.060994f
C1599 avss.n327 dvss 0.01738f
C1600 avss.n328 dvss 0.07292f
C1601 avss.n329 dvss 0.07292f
C1602 avss.n330 dvss 0.079912f
C1603 avss.n331 dvss 0.060862f
C1604 avss.t68 dvss 0.979724f
C1605 avss.n332 dvss 0.060862f
C1606 avss.n333 dvss 0.065526f
C1607 avss.n334 dvss 0.082161f
C1608 avss.n335 dvss 0.057416f
C1609 avss.n336 dvss 0.040955f
C1610 avss.n337 dvss 0.174138f
C1611 avss.n338 dvss 1.5376f
C1612 avss.n339 dvss 1.09381f
C1613 avss.n340 dvss 1.77053f
C1614 avss.n341 dvss 6.282721f
C1615 avss.n342 dvss 0.217045f
C1616 avss.n343 dvss 0.132415f
C1617 avss.n344 dvss 0.114879f
C1618 avss.n345 dvss 0.160784f
C1619 avss.n346 dvss 0.060994f
C1620 avss.n347 dvss 0.979724f
C1621 avss.t110 dvss 1.47549f
C1622 avss.t127 dvss 1.95945f
C1623 avss.t45 dvss 1.95945f
C1624 avss.t2 dvss 2.036f
C1625 avss.n348 dvss 2.44507f
C1626 avss.n349 dvss 1.08927f
C1627 avss.n350 dvss 0.783766f
C1628 avss.n351 dvss 1.73447f
.ends

