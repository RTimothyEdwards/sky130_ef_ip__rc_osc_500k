* NGSPICE file created from sky130_ef_ip__rc_osc_500k.ext - technology: sky130A

.subckt sky130_ef_ip__rc_osc_500k dout ena dvss dvdd avdd avss
X0 a_1178_9768# a_1344_7168# avss.t81 sky130_fd_pr__res_xhigh_po_0p35 l=11
X1 a_10660_3118# a_10494_518# avss.t152 sky130_fd_pr__res_xhigh_po_0p35 l=11
X2 a_4352_3118# a_4186_518# avss.t144 sky130_fd_pr__res_xhigh_po_0p35 l=11
X3 a_6490_9768# a_6656_7168# avss.t140 sky130_fd_pr__res_xhigh_po_0p35 l=11
X4 a_3502_9768# a_3336_7168# avss.t32 sky130_fd_pr__res_xhigh_po_0p35 l=11
X5 a_5162_9768# a_4996_7168# avss.t50 sky130_fd_pr__res_xhigh_po_0p35 l=11
X6 a_8814_9768# a_8648_7168# avss.t78 sky130_fd_pr__res_xhigh_po_0p35 l=11
X7 a_2692_3118# a_2858_518# avss.t73 sky130_fd_pr__res_xhigh_po_0p35 l=11
X8 a_7718_4786# ena.t0 a_7560_4786# avss.t98 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X9 a_7154_9768# a_7320_7168# avss.t97 sky130_fd_pr__res_xhigh_po_0p35 l=11
X10 a_5348_3118# a_5182_518# avss.t153 sky130_fd_pr__res_xhigh_po_0p35 l=11
X11 a_11636_7168# a_11490_518# avss.t58 sky130_fd_pr__res_xhigh_po_0p35 l=11
X12 a_4166_9768# a_4000_7168# avss.t22 sky130_fd_pr__res_xhigh_po_0p35 l=11
X13 a_11138_9768# a_11304_7168# avss.t154 sky130_fd_pr__res_xhigh_po_0p35 l=11
X14 a_4194_4788# a_3638_4788# a_4036_4788# avss.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X15 a_3688_3118# a_3854_518# avss.t24 sky130_fd_pr__res_xhigh_po_0p35 l=11
X16 a_2506_9768# a_2340_7168# avss.t94 sky130_fd_pr__res_xhigh_po_0p35 l=11
X17 a_9478_9768# a_9312_7168# avss.t108 sky130_fd_pr__res_xhigh_po_0p35 l=11
X18 a_7818_9768# a_7652_7168# avss.t76 sky130_fd_pr__res_xhigh_po_0p35 l=11
X19 a_6344_3118# a_6178_518# avss.t63 sky130_fd_pr__res_xhigh_po_0p35 l=11
X20 avdd.t15 a_2368_4788# a_2368_4788# avdd.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X21 a_1032_3118# a_866_518# avss.t23 sky130_fd_pr__res_xhigh_po_0p35 l=11
X22 a_846_9768# a_1012_7168# avss.t53 sky130_fd_pr__res_xhigh_po_0p35 l=11
X23 a_6158_9768# a_6324_7168# avss.t107 sky130_fd_pr__res_xhigh_po_0p35 l=11
X24 a_4684_3118# a_4850_518# avss.t43 sky130_fd_pr__res_xhigh_po_0p35 l=11
X25 a_10806_9768# a_10972_7168# avss.t68 sky130_fd_pr__res_xhigh_po_0p35 l=11
X26 avss.t100 ena.t1 level_shifter_0.outb_h avss.t99 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X27 a_10142_9768# a_10308_7168# avss.t25 sky130_fd_pr__res_xhigh_po_0p35 l=11
X28 a_7340_3118# a_7174_518# avss.t20 sky130_fd_pr__res_xhigh_po_0p35 l=11
X29 avdd.t13 a_2368_4788# a_4854_5653# avdd.t12 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X30 a_5826_9768# a_5992_7168# avss.t79 sky130_fd_pr__res_xhigh_po_0p35 l=11
X31 a_5162_9768# a_5328_7168# avss.t82 sky130_fd_pr__res_xhigh_po_0p35 l=11
X32 avdd.t11 a_2368_4788# a_5470_5653# avdd.t10 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X33 a_2028_3118# a_1862_518# avss.t47 sky130_fd_pr__res_xhigh_po_0p35 l=11
X34 a_5680_3118# a_5846_518# avss.t84 sky130_fd_pr__res_xhigh_po_0p35 l=11
X35 a_9146_9768# a_8980_7168# avss.t141 sky130_fd_pr__res_xhigh_po_0p35 l=11
X36 a_8336_3118# a_8170_518# avss.t35 sky130_fd_pr__res_xhigh_po_0p35 l=11
X37 a_4830_9768# a_4996_7168# avss.t60 sky130_fd_pr__res_xhigh_po_0p35 l=11
X38 a_3024_3118# a_2858_518# avss.t83 sky130_fd_pr__res_xhigh_po_0p35 l=11
X39 a_6676_3118# a_6842_518# avss.t1 sky130_fd_pr__res_xhigh_po_0p35 l=11
X40 a_1364_3118# a_1530_518# avss.t114 sky130_fd_pr__res_xhigh_po_0p35 l=11
X41 a_10474_9768# a_10640_7168# avss.t49 sky130_fd_pr__res_xhigh_po_0p35 l=11
X42 a_1842_9768# a_1676_7168# avss.t89 sky130_fd_pr__res_xhigh_po_0p35 l=11
X43 a_9332_3118# a_9166_518# avss.t27 sky130_fd_pr__res_xhigh_po_0p35 l=11
X44 a_4020_3118# a_3854_518# avss.t77 sky130_fd_pr__res_xhigh_po_0p35 l=11
X45 avdd.t22 level_shifter_0.out_h a_2368_4788# avdd.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X46 a_3082_4788# avss.t44 sky130_fd_pr__cap_mim_m3_1 l=6 w=3
X47 dvdd.t6 ena.t2 level_shifter_0.inb_l dvdd.t5 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X48 a_5494_9768# a_5660_7168# avss.t163 sky130_fd_pr__res_xhigh_po_0p35 l=11
X49 a_4750_4788# a_4194_4788# a_4854_5653# avdd.t12 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X50 a_10328_3118# a_10162_518# avss.t113 sky130_fd_pr__res_xhigh_po_0p35 l=11
X51 a_7672_3118# a_7838_518# avss.t80 sky130_fd_pr__res_xhigh_po_0p35 l=11
X52 a_1414_4786# level_shifter_0.outb_h avss.t30 avss.t29 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X53 a_4750_4788# avss.t110 sky130_fd_pr__cap_mim_m3_1 l=6 w=3
X54 a_700_3118# a_534_518# avss.t62 sky130_fd_pr__res_xhigh_po_0p35 l=11
X55 a_2360_3118# a_2526_518# avss.t0 sky130_fd_pr__res_xhigh_po_0p35 l=11
X56 a_1414_4786# level_shifter_0.out_h a_514_7168# avss.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X57 a_1032_3118# a_1198_518# avss.t115 sky130_fd_pr__res_xhigh_po_0p35 l=11
X58 a_3638_4788# avss.t36 sky130_fd_pr__cap_mim_m3_1 l=6 w=3
X59 a_5306_4788# a_4750_4788# a_5470_5653# avdd.t10 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X60 a_11324_3118# a_11158_518# avss.t95 sky130_fd_pr__res_xhigh_po_0p35 l=11
X61 a_5016_3118# a_4850_518# avss.t54 sky130_fd_pr__res_xhigh_po_0p35 l=11
X62 a_4498_9768# a_4664_7168# avss.t46 sky130_fd_pr__res_xhigh_po_0p35 l=11
X63 a_8668_3118# a_8834_518# avss.t70 sky130_fd_pr__res_xhigh_po_0p35 l=11
X64 a_9810_9768# a_9976_7168# avss.t105 sky130_fd_pr__res_xhigh_po_0p35 l=11
X65 avdd.t9 a_2368_4788# a_3622_5653# avdd.t8 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X66 a_3356_3118# a_3522_518# avss.t66 sky130_fd_pr__res_xhigh_po_0p35 l=11
X67 a_2028_3118# a_2194_518# avss.t51 sky130_fd_pr__res_xhigh_po_0p35 l=11
X68 a_6260_4788# a_1414_4786# avss.t19 avss.t18 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X69 a_5306_4788# avss.t164 sky130_fd_pr__cap_mim_m3_1 l=6 w=3
X70 a_3170_9768# a_3004_7168# avss.t160 sky130_fd_pr__res_xhigh_po_0p35 l=11
X71 a_6012_3118# a_5846_518# avss.t48 sky130_fd_pr__res_xhigh_po_0p35 l=11
X72 a_1510_9768# a_1344_7168# avss.t55 sky130_fd_pr__res_xhigh_po_0p35 l=11
X73 a_6822_9768# a_6656_7168# avss.t96 sky130_fd_pr__res_xhigh_po_0p35 l=11
X74 a_8482_9768# a_8316_7168# avss.t86 sky130_fd_pr__res_xhigh_po_0p35 l=11
X75 avdd.t7 a_2368_4788# a_3006_5653# avdd.t6 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X76 a_9664_3118# a_9830_518# avss.t165 sky130_fd_pr__res_xhigh_po_0p35 l=11
X77 avdd.t5 a_2368_4788# a_4238_5653# avdd.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X78 dvss.t7 ena.t3 level_shifter_0.inb_l dvss.t6 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X79 a_10806_9768# a_10640_7168# avss.t57 sky130_fd_pr__res_xhigh_po_0p35 l=11
X80 a_9482_5327# level_shifter_0.out_h level_shifter_0.outb_h avdd.t21 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X81 a_3024_3118# a_3190_518# avss.t166 sky130_fd_pr__res_xhigh_po_0p35 l=11
X82 a_3502_9768# a_3668_7168# avss.t106 sky130_fd_pr__res_xhigh_po_0p35 l=11
X83 avdd.t3 a_2368_4788# a_6702_5653# avdd.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X84 a_4352_3118# a_4518_518# avss.t109 sky130_fd_pr__res_xhigh_po_0p35 l=11
X85 a_2174_9768# a_2008_7168# avss.t52 sky130_fd_pr__res_xhigh_po_0p35 l=11
X86 a_7486_9768# a_7320_7168# avss.t150 sky130_fd_pr__res_xhigh_po_0p35 l=11
X87 a_10660_3118# a_10826_518# avss.t121 sky130_fd_pr__res_xhigh_po_0p35 l=11
X88 a_5826_9768# a_5660_7168# avss.t126 sky130_fd_pr__res_xhigh_po_0p35 l=11
X89 dout.t1 a_7718_4786# dvdd.t1 dvdd.t0 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X90 a_7008_3118# a_6842_518# avss.t127 sky130_fd_pr__res_xhigh_po_0p35 l=11
X91 a_1696_3118# a_1530_518# avss.t122 sky130_fd_pr__res_xhigh_po_0p35 l=11
X92 avdd.t1 a_2368_4788# a_6086_5653# avdd.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X93 a_9332_3118# a_9498_518# avss.t130 sky130_fd_pr__res_xhigh_po_0p35 l=11
X94 a_11890_5939# a_7718_4786# dvss.t3 dvss.t2 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.15
D0 dvss.t5 ena.t4 sky130_fd_pr__diode_pw2nd_05v5 pj=1.8e+06 area=2.025e+11
X95 a_4166_9768# a_4332_7168# avss.t117 sky130_fd_pr__res_xhigh_po_0p35 l=11
X96 a_5348_3118# a_5514_518# avss.t119 sky130_fd_pr__res_xhigh_po_0p35 l=11
X97 a_4020_3118# a_4186_518# avss.t120 sky130_fd_pr__res_xhigh_po_0p35 l=11
X98 a_9478_9768# a_9644_7168# avss.t116 sky130_fd_pr__res_xhigh_po_0p35 l=11
X99 a_10328_3118# a_10494_518# avss.t129 sky130_fd_pr__res_xhigh_po_0p35 l=11
X100 a_514_9768# a_680_7168# avss.t136 sky130_fd_pr__res_xhigh_po_0p35 l=11
X101 level_shifter_0.out_h level_shifter_0.outb_h a_8714_4659# avdd.t18 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X102 a_1178_9768# a_1012_7168# avss.t135 sky130_fd_pr__res_xhigh_po_0p35 l=11
X103 a_8004_3118# a_7838_518# avss.t138 sky130_fd_pr__res_xhigh_po_0p35 l=11
X104 a_2692_3118# a_2526_518# avss.t128 sky130_fd_pr__res_xhigh_po_0p35 l=11
X105 a_5148_4788# a_1414_4786# avss.t17 avss.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X106 a_2982_4700# a_5862_4788# a_6260_4788# avss.t18 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X107 a_8150_9768# a_7984_7168# avss.t134 sky130_fd_pr__res_xhigh_po_0p35 l=11
X108 level_shifter_0.out_h level_shifter_0.inb_l avss.t75 avss.t74 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X109 a_5704_4788# a_1414_4786# avss.t15 avss.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X110 a_6344_3118# a_6510_518# avss.t149 sky130_fd_pr__res_xhigh_po_0p35 l=11
X111 a_3638_4788# a_3082_4788# a_3622_5653# avdd.t8 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X112 a_11324_3118# a_11490_518# avss.t137 sky130_fd_pr__res_xhigh_po_0p35 l=11
X113 a_5016_3118# a_5182_518# avss.t142 sky130_fd_pr__res_xhigh_po_0p35 l=11
X114 a_700_3118# a_866_518# avss.t125 sky130_fd_pr__res_xhigh_po_0p35 l=11
X115 a_9000_3118# a_8834_518# avss.t124 sky130_fd_pr__res_xhigh_po_0p35 l=11
X116 dvss.t1 level_shifter_0.inb_l dout.t0 dvss.t0 sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.15
X117 a_3480_4788# a_1414_4786# avss.t13 avss.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X118 a_3170_9768# a_3336_7168# avss.t143 sky130_fd_pr__res_xhigh_po_0p35 l=11
X119 a_8482_9768# a_8648_7168# avss.t118 sky130_fd_pr__res_xhigh_po_0p35 l=11
X120 a_3082_4788# a_2982_4700# a_3006_5653# avdd.t6 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X121 a_4194_4788# a_3638_4788# a_4238_5653# avdd.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X122 dvdd.t4 ena.t5 a_7718_4786# dvdd.t3 sky130_fd_pr__pfet_01v8 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.15
X123 a_7154_9768# a_6988_7168# avss.t146 sky130_fd_pr__res_xhigh_po_0p35 l=11
X124 a_3688_3118# a_3522_518# avss.t123 sky130_fd_pr__res_xhigh_po_0p35 l=11
X125 a_11138_9768# a_10972_7168# avss.t148 sky130_fd_pr__res_xhigh_po_0p35 l=11
X126 a_2982_4700# a_5862_4788# a_6702_5653# avdd.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X127 a_7340_3118# a_7506_518# avss.t90 sky130_fd_pr__res_xhigh_po_0p35 l=11
X128 a_6012_3118# a_6178_518# avss.t41 sky130_fd_pr__res_xhigh_po_0p35 l=11
X129 a_3834_9768# a_4000_7168# avss.t64 sky130_fd_pr__res_xhigh_po_0p35 l=11
X130 a_9146_9768# a_9312_7168# avss.t157 sky130_fd_pr__res_xhigh_po_0p35 l=11
X131 a_9996_3118# a_9830_518# avss.t69 sky130_fd_pr__res_xhigh_po_0p35 l=11
X132 a_4684_3118# a_4518_518# avss.t147 sky130_fd_pr__res_xhigh_po_0p35 l=11
X133 a_5862_4788# a_5306_4788# a_6086_5653# avdd.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X134 a_10992_3118# a_10826_518# avss.t93 sky130_fd_pr__res_xhigh_po_0p35 l=11
X135 a_8336_3118# a_8502_518# avss.t67 sky130_fd_pr__res_xhigh_po_0p35 l=11
X136 a_6158_9768# a_5992_7168# avss.t101 sky130_fd_pr__res_xhigh_po_0p35 l=11
X137 a_5306_4788# a_4750_4788# a_5148_4788# avss.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X138 a_7008_3118# a_7174_518# avss.t56 sky130_fd_pr__res_xhigh_po_0p35 l=11
X139 a_7718_4786# a_2982_4700# dvdd.t2 avdd.t23 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X140 a_4592_4788# a_1414_4786# avss.t11 avss.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X141 a_5862_4788# a_5306_4788# a_5704_4788# avss.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X142 a_846_9768# a_680_7168# avss.t65 sky130_fd_pr__res_xhigh_po_0p35 l=11
X143 a_8814_9768# a_8980_7168# avss.t112 sky130_fd_pr__res_xhigh_po_0p35 l=11
X144 a_5680_3118# a_5514_518# avss.t85 sky130_fd_pr__res_xhigh_po_0p35 l=11
X145 a_2838_9768# a_3004_7168# avss.t102 sky130_fd_pr__res_xhigh_po_0p35 l=11
X146 avdd.t20 level_shifter_0.out_h a_8714_4659# avdd.t18 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X147 a_8150_9768# a_8316_7168# avss.t139 sky130_fd_pr__res_xhigh_po_0p35 l=11
X148 a_3638_4788# a_3082_4788# a_3480_4788# avss.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X149 a_2526_4188# a_1414_4786# avss.t9 avss.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X150 a_8004_3118# a_8170_518# avss.t39 sky130_fd_pr__res_xhigh_po_0p35 l=11
X151 a_2924_4788# a_1414_4786# avss.t7 avss.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X152 a_11470_9768# a_11304_7168# avss.t159 sky130_fd_pr__res_xhigh_po_0p35 l=11
X153 a_9482_5327# level_shifter_0.outb_h avdd.t17 avdd.t16 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X154 a_2506_9768# a_2672_7168# avss.t40 sky130_fd_pr__res_xhigh_po_0p35 l=11
X155 a_7818_9768# a_7984_7168# avss.t145 sky130_fd_pr__res_xhigh_po_0p35 l=11
X156 a_11890_5939# ena.t6 dout.t2 dvss.t4 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.15
X157 a_1842_9768# a_2008_7168# avss.t155 sky130_fd_pr__res_xhigh_po_0p35 l=11
X158 a_6676_3118# a_6510_518# avss.t161 sky130_fd_pr__res_xhigh_po_0p35 l=11
X159 a_6490_9768# a_6324_7168# avss.t72 sky130_fd_pr__res_xhigh_po_0p35 l=11
X160 a_1364_3118# a_1198_518# avss.t162 sky130_fd_pr__res_xhigh_po_0p35 l=11
X161 a_4830_9768# a_4664_7168# avss.t45 sky130_fd_pr__res_xhigh_po_0p35 l=11
X162 a_9000_3118# a_9166_518# avss.t156 sky130_fd_pr__res_xhigh_po_0p35 l=11
X163 a_10474_9768# a_10308_7168# avss.t92 sky130_fd_pr__res_xhigh_po_0p35 l=11
X164 a_9996_3118# a_10162_518# avss.t133 sky130_fd_pr__res_xhigh_po_0p35 l=11
X165 a_1510_9768# a_1676_7168# avss.t28 sky130_fd_pr__res_xhigh_po_0p35 l=11
X166 a_7672_3118# a_7506_518# avss.t132 sky130_fd_pr__res_xhigh_po_0p35 l=11
X167 a_514_9768# a_514_7168# avss.t21 sky130_fd_pr__res_xhigh_po_0p35 l=11
X168 a_6822_9768# a_6988_7168# avss.t34 sky130_fd_pr__res_xhigh_po_0p35 l=11
X169 a_4750_4788# a_4194_4788# a_4592_4788# avss.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X170 a_2360_3118# a_2194_518# avss.t103 sky130_fd_pr__res_xhigh_po_0p35 l=11
X171 a_4194_4788# avss.t31 sky130_fd_pr__cap_mim_m3_1 l=6 w=3
X172 a_5494_9768# a_5328_7168# avss.t33 sky130_fd_pr__res_xhigh_po_0p35 l=11
X173 a_2526_4188# level_shifter_0.out_h a_2368_4788# avss.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X174 a_3834_9768# a_3668_7168# avss.t88 sky130_fd_pr__res_xhigh_po_0p35 l=11
X175 a_3082_4788# a_2982_4700# a_2924_4788# avss.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X176 avdd a_534_518# avss.t38 sky130_fd_pr__res_xhigh_po_0p35 l=11
X177 a_1414_4786# a_1414_4786# avss.t5 avss.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X178 a_7560_4786# a_2982_4700# avss.t131 avss.t98 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X179 a_2174_9768# a_2340_7168# avss.t71 sky130_fd_pr__res_xhigh_po_0p35 l=11
X180 a_7486_9768# a_7652_7168# avss.t26 sky130_fd_pr__res_xhigh_po_0p35 l=11
X181 a_10992_3118# a_11158_518# avss.t158 sky130_fd_pr__res_xhigh_po_0p35 l=11
X182 a_8668_3118# a_8502_518# avss.t151 sky130_fd_pr__res_xhigh_po_0p35 l=11
X183 a_3356_3118# a_3190_518# avss.t61 sky130_fd_pr__res_xhigh_po_0p35 l=11
X184 a_4036_4788# a_1414_4786# avss.t3 avss.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X185 a_11470_9768# a_11636_7168# avss.t111 sky130_fd_pr__res_xhigh_po_0p35 l=11
X186 a_2838_9768# a_2672_7168# avss.t37 sky130_fd_pr__res_xhigh_po_0p35 l=11
X187 a_4498_9768# a_4332_7168# avss.t87 sky130_fd_pr__res_xhigh_po_0p35 l=11
X188 a_9810_9768# a_9644_7168# avss.t91 sky130_fd_pr__res_xhigh_po_0p35 l=11
X189 a_1696_3118# a_1862_518# avss.t59 sky130_fd_pr__res_xhigh_po_0p35 l=11
X190 a_9664_3118# a_9498_518# avss.t104 sky130_fd_pr__res_xhigh_po_0p35 l=11
X191 a_10142_9768# a_9976_7168# avss.t42 sky130_fd_pr__res_xhigh_po_0p35 l=11
R0 avss.n269 avss.n3 49093.8
R1 avss.n348 avss.n3 49093.8
R2 avss.n348 avss.n4 49093.8
R3 avss.n269 avss.n4 49093.8
R4 avss.n36 avss.n28 49093.8
R5 avss.n322 avss.n28 49093.8
R6 avss.n322 avss.n29 49093.8
R7 avss.n36 avss.n29 49093.8
R8 avss.n300 avss.n299 4540.48
R9 avss.n324 avss.n323 3194
R10 avss.n301 avss.n39 1647.1
R11 avss.n301 avss.n40 1647.1
R12 avss.n314 avss.n40 1647.1
R13 avss.n314 avss.n39 1647.1
R14 avss.n346 avss.n5 1647.1
R15 avss.n346 avss.n6 1647.1
R16 avss.n326 avss.n6 1647.1
R17 avss.n326 avss.n5 1647.1
R18 avss.n331 avss.n22 1647.1
R19 avss.n332 avss.n22 1647.1
R20 avss.n332 avss.n21 1647.1
R21 avss.n331 avss.n21 1647.1
R22 avss.n215 avss.n214 1647.1
R23 avss.n220 avss.n215 1647.1
R24 avss.n221 avss.n220 1647.1
R25 avss.n221 avss.n214 1647.1
R26 avss.n235 avss.n105 1647.1
R27 avss.n234 avss.n105 1647.1
R28 avss.n234 avss.n104 1647.1
R29 avss.n235 avss.n104 1647.1
R30 avss.n240 avss.n98 1647.1
R31 avss.n241 avss.n98 1647.1
R32 avss.n241 avss.n97 1647.1
R33 avss.n240 avss.n97 1647.1
R34 avss.n189 avss.n182 1647.1
R35 avss.n182 avss.n123 1647.1
R36 avss.n178 avss.n123 1647.1
R37 avss.n189 avss.n178 1647.1
R38 avss.n253 avss.n81 1647.1
R39 avss.n252 avss.n81 1647.1
R40 avss.n252 avss.n80 1647.1
R41 avss.n253 avss.n80 1647.1
R42 avss.n258 avss.n74 1647.1
R43 avss.n259 avss.n74 1647.1
R44 avss.n259 avss.n73 1647.1
R45 avss.n258 avss.n73 1647.1
R46 avss.n162 avss.n140 1647.1
R47 avss.n140 avss.n135 1647.1
R48 avss.n136 avss.n135 1647.1
R49 avss.n162 avss.n136 1647.1
R50 avss.n156 avss.n57 1647.1
R51 avss.n156 avss.n58 1647.1
R52 avss.n288 avss.n58 1647.1
R53 avss.n288 avss.n57 1647.1
R54 avss.n290 avss.n49 1647.1
R55 avss.n290 avss.n50 1647.1
R56 avss.n297 avss.n50 1647.1
R57 avss.n297 avss.n49 1647.1
R58 avss.n202 avss.n18 1647.1
R59 avss.n202 avss.n23 1647.1
R60 avss.n217 avss.n23 1647.1
R61 avss.n217 avss.n18 1647.1
R62 avss.n216 avss.n200 1647.1
R63 avss.n216 avss.n208 1647.1
R64 avss.n223 avss.n208 1647.1
R65 avss.n223 avss.n200 1647.1
R66 avss.n209 avss.n106 1647.1
R67 avss.n209 avss.n107 1647.1
R68 avss.n114 avss.n107 1647.1
R69 avss.n114 avss.n106 1647.1
R70 avss.n117 avss.n95 1647.1
R71 avss.n117 avss.n99 1647.1
R72 avss.n179 avss.n99 1647.1
R73 avss.n179 avss.n95 1647.1
R74 avss.n122 avss.n121 1647.1
R75 avss.n190 avss.n121 1647.1
R76 avss.n190 avss.n120 1647.1
R77 avss.n122 avss.n120 1647.1
R78 avss.n175 avss.n82 1647.1
R79 avss.n175 avss.n83 1647.1
R80 avss.n126 avss.n83 1647.1
R81 avss.n126 avss.n82 1647.1
R82 avss.n129 avss.n71 1647.1
R83 avss.n129 avss.n75 1647.1
R84 avss.n137 avss.n75 1647.1
R85 avss.n137 avss.n71 1647.1
R86 avss.n134 avss.n133 1647.1
R87 avss.n163 avss.n133 1647.1
R88 avss.n163 avss.n132 1647.1
R89 avss.n134 avss.n132 1647.1
R90 avss.n152 avss.n62 1647.1
R91 avss.n152 avss.n144 1647.1
R92 avss.n144 avss.n56 1647.1
R93 avss.n62 avss.n56 1647.1
R94 avss.n292 avss.n54 1647.1
R95 avss.n55 avss.n54 1647.1
R96 avss.n55 avss.n48 1647.1
R97 avss.n292 avss.n48 1647.1
R98 avss.n308 avss.n45 1647.1
R99 avss.n310 avss.n44 1647.1
R100 avss.n310 avss.n45 1647.1
R101 avss.n321 avss.n30 1079.34
R102 avss.n270 avss.n2 1068.09
R103 avss.n349 avss.n2 1063.11
R104 avss.n31 avss.n30 1048.5
R105 avss.t99 avss.n35 934.398
R106 avss.n300 avss.t74 934.398
R107 avss.n321 avss.n320 917.9
R108 avss.n271 avss.n268 883.951
R109 avss.n315 avss.n38 697.509
R110 avss.n309 avss.n44 613.538
R111 avss.n319 avss.n31 612.216
R112 avss.n316 avss.n35 552.742
R113 avss.n350 avss.n1 479.428
R114 avss.n320 avss.n319 434.247
R115 avss.n267 avss.n1 408.832
R116 avss.n64 avss.t131 348.699
R117 avss.n343 avss.t30 347.341
R118 avss.n283 avss.t19 346.911
R119 avss.n264 avss.t15 346.911
R120 avss.n87 avss.t17 346.911
R121 avss.n249 avss.t11 346.911
R122 avss.n246 avss.t3 346.911
R123 avss.n227 avss.t13 346.911
R124 avss.n231 avss.t7 346.911
R125 avss.n337 avss.t9 346.911
R126 avss.n19 avss.t5 346.889
R127 avss.n46 avss.t100 346.827
R128 avss.n33 avss.t75 346.815
R129 avss.n316 avss.n315 236.889
R130 avss.t74 avss.n38 236.889
R131 avss.t58 avss.t137 213.194
R132 avss.t137 avss.t95 213.194
R133 avss.t95 avss.t158 213.194
R134 avss.t158 avss.t93 213.194
R135 avss.t93 avss.t121 213.194
R136 avss.t121 avss.t152 213.194
R137 avss.t152 avss.t129 213.194
R138 avss.t129 avss.t113 213.194
R139 avss.t113 avss.t133 213.194
R140 avss.t133 avss.t69 213.194
R141 avss.t69 avss.t165 213.194
R142 avss.t159 avss.t111 212.946
R143 avss.t154 avss.t159 212.946
R144 avss.t148 avss.t154 212.946
R145 avss.t68 avss.t148 212.946
R146 avss.t57 avss.t68 212.946
R147 avss.t49 avss.t57 212.946
R148 avss.t92 avss.t49 212.946
R149 avss.t25 avss.t92 212.946
R150 avss.t42 avss.t25 212.946
R151 avss.t105 avss.t42 212.946
R152 avss.t91 avss.t105 212.946
R153 avss.n293 avss.n292 210
R154 avss.n292 avss.t98 210
R155 avss.n146 avss.n55 210
R156 avss.t98 avss.n55 210
R157 avss.n285 avss.n62 210
R158 avss.t18 avss.n62 210
R159 avss.n149 avss.n144 210
R160 avss.n144 avss.t18 210
R161 avss.n134 avss.n66 210
R162 avss.t14 avss.n134 210
R163 avss.n164 avss.n163 210
R164 avss.n163 avss.t14 210
R165 avss.n260 avss.n71 210
R166 avss.t16 avss.n71 210
R167 avss.n167 avss.n75 210
R168 avss.t16 avss.n75 210
R169 avss.n251 avss.n82 210
R170 avss.t10 avss.n82 210
R171 avss.n170 avss.n83 210
R172 avss.t10 avss.n83 210
R173 avss.n122 avss.n90 210
R174 avss.t2 avss.n122 210
R175 avss.n191 avss.n190 210
R176 avss.n190 avss.t2 210
R177 avss.n242 avss.n95 210
R178 avss.t12 avss.n95 210
R179 avss.n194 avss.n99 210
R180 avss.t12 avss.n99 210
R181 avss.n233 avss.n106 210
R182 avss.t6 avss.n106 210
R183 avss.n197 avss.n107 210
R184 avss.t6 avss.n107 210
R185 avss.n200 avss.n13 210
R186 avss.t8 avss.n200 210
R187 avss.n208 avss.n207 210
R188 avss.t8 avss.n208 210
R189 avss.n333 avss.n18 210
R190 avss.t4 avss.n18 210
R191 avss.n204 avss.n23 210
R192 avss.t4 avss.n23 210
R193 avss.n295 avss.n49 210
R194 avss.t98 avss.n49 210
R195 avss.n293 avss.n50 210
R196 avss.t98 avss.n50 210
R197 avss.n61 avss.n57 210
R198 avss.t18 avss.n57 210
R199 avss.n285 avss.n58 210
R200 avss.t18 avss.n58 210
R201 avss.n162 avss.n161 210
R202 avss.t14 avss.n162 210
R203 avss.n135 avss.n66 210
R204 avss.t14 avss.n135 210
R205 avss.n258 avss.n257 210
R206 avss.t16 avss.n258 210
R207 avss.n260 avss.n259 210
R208 avss.n259 avss.t16 210
R209 avss.n254 avss.n253 210
R210 avss.n253 avss.t10 210
R211 avss.n252 avss.n251 210
R212 avss.t10 avss.n252 210
R213 avss.n189 avss.n188 210
R214 avss.t2 avss.n189 210
R215 avss.n123 avss.n90 210
R216 avss.t2 avss.n123 210
R217 avss.n240 avss.n239 210
R218 avss.t12 avss.n240 210
R219 avss.n242 avss.n241 210
R220 avss.n241 avss.t12 210
R221 avss.n236 avss.n235 210
R222 avss.n235 avss.t6 210
R223 avss.n234 avss.n233 210
R224 avss.t6 avss.n234 210
R225 avss.n214 avss.n213 210
R226 avss.t8 avss.n214 210
R227 avss.n220 avss.n13 210
R228 avss.n220 avss.t8 210
R229 avss.n331 avss.n330 210
R230 avss.t4 avss.n331 210
R231 avss.n333 avss.n332 210
R232 avss.n332 avss.t4 210
R233 avss.n7 avss.n5 210
R234 avss.t29 avss.n5 210
R235 avss.n8 avss.n6 210
R236 avss.t29 avss.n6 210
R237 avss.n304 avss.n39 210
R238 avss.t74 avss.n39 210
R239 avss.n42 avss.n40 210
R240 avss.t74 avss.n40 210
R241 avss.n311 avss.n310 210
R242 avss.n310 avss.t99 210
R243 avss.n308 avss.n307 210
R244 avss.n269 avss.t58 208.338
R245 avss.t111 avss.n36 208.115
R246 avss.t116 avss.t91 204.929
R247 avss.t165 avss.t104 204.137
R248 avss.t108 avss.t116 197.994
R249 avss.t157 avss.t108 197.994
R250 avss.t141 avss.t157 197.994
R251 avss.t112 avss.t141 197.994
R252 avss.t78 avss.t118 197.994
R253 avss.t118 avss.t86 197.994
R254 avss.t86 avss.t139 197.994
R255 avss.t139 avss.t134 197.994
R256 avss.t134 avss.t145 197.994
R257 avss.t145 avss.t76 197.994
R258 avss.t76 avss.t26 197.994
R259 avss.t26 avss.t150 197.994
R260 avss.t150 avss.t97 197.994
R261 avss.t97 avss.t146 197.994
R262 avss.t146 avss.t34 197.964
R263 avss.t34 avss.t96 197.94
R264 avss.t96 avss.t140 197.94
R265 avss.t140 avss.t72 197.94
R266 avss.t72 avss.t107 197.94
R267 avss.t107 avss.t101 197.94
R268 avss.t79 avss.t126 197.94
R269 avss.t126 avss.t163 197.94
R270 avss.t163 avss.t33 197.94
R271 avss.t33 avss.t82 197.94
R272 avss.t82 avss.t50 197.94
R273 avss.t50 avss.t60 197.94
R274 avss.t60 avss.t45 197.94
R275 avss.t45 avss.t46 197.94
R276 avss.t46 avss.t87 197.94
R277 avss.t87 avss.t117 197.94
R278 avss.t117 avss.t22 197.94
R279 avss.t22 avss.t64 197.94
R280 avss.t64 avss.t88 197.94
R281 avss.t88 avss.t106 197.94
R282 avss.t106 avss.t32 197.94
R283 avss.t32 avss.t143 197.94
R284 avss.t143 avss.t160 197.94
R285 avss.t160 avss.t102 197.94
R286 avss.t102 avss.t37 197.94
R287 avss.t37 avss.t40 197.94
R288 avss.t40 avss.t94 197.94
R289 avss.t94 avss.t71 197.94
R290 avss.t71 avss.t52 197.94
R291 avss.t52 avss.t155 197.94
R292 avss.t155 avss.t89 197.94
R293 avss.t89 avss.t28 197.94
R294 avss.t28 avss.t55 197.94
R295 avss.t55 avss.t81 197.94
R296 avss.t135 avss.t53 197.94
R297 avss.t53 avss.t65 197.94
R298 avss.t65 avss.t136 197.94
R299 avss.t136 avss.t21 197.94
R300 avss.t21 avss.n322 194.738
R301 avss.t104 avss.t130 191.405
R302 avss.t130 avss.t27 191.405
R303 avss.t27 avss.t156 191.405
R304 avss.t156 avss.t124 191.405
R305 avss.t124 avss.t70 191.405
R306 avss.t70 avss.t151 191.405
R307 avss.t151 avss.t67 191.405
R308 avss.n145 avss.n48 168.274
R309 avss.n298 avss.n48 168
R310 avss.n54 avss.n52 168
R311 avss.n291 avss.n54 168
R312 avss.n59 avss.n56 168
R313 avss.n289 avss.n56 168
R314 avss.n152 avss.n151 168
R315 avss.n155 avss.n152 168
R316 avss.n141 avss.n132 168
R317 avss.n153 avss.n132 168
R318 avss.n133 avss.n68 168
R319 avss.n139 avss.n133 168
R320 avss.n137 avss.n70 168
R321 avss.n138 avss.n137 168
R322 avss.n130 avss.n129 168
R323 avss.n129 avss.n128 168
R324 avss.n126 avss.n124 168
R325 avss.n127 avss.n126 168
R326 avss.n175 avss.n174 168
R327 avss.n176 avss.n175 168
R328 avss.n183 avss.n120 168
R329 avss.n177 avss.n120 168
R330 avss.n121 avss.n92 168
R331 avss.n181 avss.n121 168
R332 avss.n179 avss.n94 168
R333 avss.n180 avss.n179 168
R334 avss.n118 avss.n117 168
R335 avss.n117 avss.n116 168
R336 avss.n114 avss.n112 168
R337 avss.n115 avss.n114 168
R338 avss.n209 avss.n110 168
R339 avss.n210 avss.n209 168
R340 avss.n224 avss.n223 168
R341 avss.n223 avss.n222 168
R342 avss.n216 avss.n15 168
R343 avss.n219 avss.n216 168
R344 avss.n217 avss.n17 168
R345 avss.n218 avss.n217 168
R346 avss.n203 avss.n202 168
R347 avss.n202 avss.n27 168
R348 avss.n297 avss.n296 168
R349 avss.n298 avss.n297 168
R350 avss.n290 avss.n53 168
R351 avss.n291 avss.n290 168
R352 avss.n288 avss.n287 168
R353 avss.n289 avss.n288 168
R354 avss.n157 avss.n156 168
R355 avss.n156 avss.n155 168
R356 avss.n143 avss.n136 168
R357 avss.n153 avss.n136 168
R358 avss.n140 avss.n67 168
R359 avss.n140 avss.n139 168
R360 avss.n73 avss.n69 168
R361 avss.n138 avss.n73 168
R362 avss.n77 avss.n74 168
R363 avss.n128 avss.n74 168
R364 avss.n80 avss.n78 168
R365 avss.n127 avss.n80 168
R366 avss.n85 avss.n81 168
R367 avss.n176 avss.n81 168
R368 avss.n185 avss.n178 168
R369 avss.n178 avss.n177 168
R370 avss.n182 avss.n91 168
R371 avss.n182 avss.n181 168
R372 avss.n97 avss.n93 168
R373 avss.n180 avss.n97 168
R374 avss.n101 avss.n98 168
R375 avss.n116 avss.n98 168
R376 avss.n104 avss.n102 168
R377 avss.n115 avss.n104 168
R378 avss.n109 avss.n105 168
R379 avss.n210 avss.n105 168
R380 avss.n221 avss.n111 168
R381 avss.n222 avss.n221 168
R382 avss.n215 avss.n14 168
R383 avss.n219 avss.n215 168
R384 avss.n21 avss.n16 168
R385 avss.n218 avss.n21 168
R386 avss.n25 avss.n22 168
R387 avss.n27 avss.n22 168
R388 avss.n327 avss.n326 168
R389 avss.n326 avss.n325 168
R390 avss.n346 avss.n345 168
R391 avss.n347 avss.n346 168
R392 avss.n302 avss.n301 168
R393 avss.n301 avss.n300 168
R394 avss.n45 avss.n41 168
R395 avss.n45 avss.n35 168
R396 avss.n314 avss.n313 168
R397 avss.n315 avss.n314 168
R398 avss.n44 avss.n43 168
R399 avss.n38 avss.t112 163.405
R400 avss.n348 avss.t38 147.621
R401 avss.n323 avss.t81 146.667
R402 avss.t39 avss.t138 145.094
R403 avss.t132 avss.t80 145.094
R404 avss.t20 avss.t56 145.094
R405 avss.t56 avss.t127 145.094
R406 avss.t127 avss.t1 145.094
R407 avss.t1 avss.t161 145.094
R408 avss.t63 avss.t149 145.094
R409 avss.t54 avss.t142 145.094
R410 avss.t43 avss.t147 145.094
R411 avss.t61 avss.t66 145.094
R412 avss.t166 avss.t83 145.094
R413 avss.t122 avss.t59 145.094
R414 avss.t114 avss.t162 145.094
R415 avss.t125 avss.t23 145.094
R416 avss.t62 avss.t125 145.094
R417 avss.t38 avss.t62 145.094
R418 avss.t138 avss.n298 138.101
R419 avss.t67 avss.t35 136.425
R420 avss.t18 avss.t41 135.48
R421 avss.n204 avss.n203 131.274
R422 avss.t10 avss.t109 128.487
R423 avss.n153 avss.t84 125.865
R424 avss.t4 avss.t47 124.99
R425 avss.t6 avss.t73 121.495
R426 avss.n177 avss.t120 118.873
R427 avss.t12 avss.t123 117.999
R428 avss.n309 avss.n308 116.876
R429 avss.t103 avss.n219 115.376
R430 avss.t161 avss.n289 113.627
R431 avss.n128 avss.n127 113.627
R432 avss.n116 avss.n115 113.627
R433 avss.n325 avss.n27 113.627
R434 avss.n222 avss.t0 111.879
R435 avss.t98 avss.t90 111.005
R436 avss.t16 avss.t153 111.005
R437 avss.n294 avss.n52 109.501
R438 avss.n287 avss.n59 109.001
R439 avss.n328 avss.n327 109.001
R440 avss.n327 avss.n26 109.001
R441 avss.n151 avss.n63 109.001
R442 avss.n225 avss.n111 109.001
R443 avss.n225 avss.n224 109.001
R444 avss.n335 avss.n14 109.001
R445 avss.n335 avss.n15 109.001
R446 avss.n108 avss.n102 109.001
R447 avss.n112 avss.n108 109.001
R448 avss.n226 avss.n109 109.001
R449 avss.n226 avss.n110 109.001
R450 avss.n243 avss.n93 109.001
R451 avss.n243 avss.n94 109.001
R452 avss.n113 avss.n101 109.001
R453 avss.n118 avss.n113 109.001
R454 avss.n185 avss.n184 109.001
R455 avss.n184 avss.n183 109.001
R456 avss.n244 avss.n91 109.001
R457 avss.n244 avss.n92 109.001
R458 avss.n84 avss.n78 109.001
R459 avss.n124 avss.n84 109.001
R460 avss.n86 avss.n85 109.001
R461 avss.n174 avss.n86 109.001
R462 avss.n261 avss.n69 109.001
R463 avss.n261 avss.n70 109.001
R464 avss.n125 avss.n77 109.001
R465 avss.n130 avss.n125 109.001
R466 avss.n143 avss.n142 109.001
R467 avss.n142 avss.n141 109.001
R468 avss.n262 avss.n67 109.001
R469 avss.n262 avss.n68 109.001
R470 avss.n157 avss.n63 109.001
R471 avss.n329 avss.n25 109.001
R472 avss.n201 avss.n25 109.001
R473 avss.n24 avss.n16 109.001
R474 avss.n334 avss.n16 109.001
R475 avss.n334 avss.n17 109.001
R476 avss.n203 avss.n201 109.001
R477 avss.n317 avss.n316 108.63
R478 avss.n148 avss.n59 108.501
R479 avss.n151 avss.n150 108.501
R480 avss.n211 avss.n111 108.501
R481 avss.n224 avss.n199 108.501
R482 avss.n212 avss.n14 108.501
R483 avss.n206 avss.n15 108.501
R484 avss.n237 avss.n102 108.501
R485 avss.n196 avss.n112 108.501
R486 avss.n109 avss.n103 108.501
R487 avss.n198 avss.n110 108.501
R488 avss.n100 avss.n93 108.501
R489 avss.n193 avss.n94 108.501
R490 avss.n238 avss.n101 108.501
R491 avss.n195 avss.n118 108.501
R492 avss.n186 avss.n185 108.501
R493 avss.n183 avss.n119 108.501
R494 avss.n187 avss.n91 108.501
R495 avss.n192 avss.n92 108.501
R496 avss.n255 avss.n78 108.501
R497 avss.n169 avss.n124 108.501
R498 avss.n85 avss.n79 108.501
R499 avss.n174 avss.n173 108.501
R500 avss.n76 avss.n69 108.501
R501 avss.n166 avss.n70 108.501
R502 avss.n256 avss.n77 108.501
R503 avss.n168 avss.n130 108.501
R504 avss.n159 avss.n143 108.501
R505 avss.n141 avss.n131 108.501
R506 avss.n160 avss.n67 108.501
R507 avss.n165 avss.n68 108.501
R508 avss.n158 avss.n157 108.501
R509 avss.n205 avss.n17 108.501
R510 avss.n181 avss.t77 108.383
R511 avss.n147 avss.n52 107.501
R512 avss.n299 avss.t35 104.888
R513 avss.n139 avss.t85 101.391
R514 avss.t101 avss.n37 98.9707
R515 avss.n37 avss.t79 98.9707
R516 avss.t29 avss.n324 94.3986
R517 avss.n148 avss.n147 93.447
R518 avss.t144 avss.n176 87.4061
R519 avss.t14 avss.t85 84.784
R520 avss.t51 avss.n218 83.9099
R521 avss.t128 avss.n210 80.4137
R522 avss.t99 avss.n309 78.2248
R523 avss.t2 avss.t77 77.7915
R524 avss.t24 avss.n180 76.9175
R525 avss.t90 avss.n291 75.1694
R526 avss.n138 avss.t153 75.1694
R527 avss.t8 avss.t0 74.2953
R528 avss.t23 avss.n347 73.4212
R529 avss.n154 avss.t48 72.5472
R530 avss.n347 avss.t115 71.6731
R531 avss.t8 avss.t103 70.7991
R532 avss.n291 avss.t20 69.925
R533 avss.t119 avss.n138 69.925
R534 avss.n180 avss.t123 68.1769
R535 avss.t2 avss.t120 67.3028
R536 avss.n311 avss.n43 66.8168
R537 avss.n302 avss.n42 66.5469
R538 avss.n210 avss.t73 64.6807
R539 avss.n218 avss.t47 61.1844
R540 avss.t14 avss.t84 60.3104
R541 avss.n176 avss.t109 57.6882
R542 avss.n296 avss.n295 57.3558
R543 avss.n345 avss.n7 54.9135
R544 avss.n303 avss.n302 53.7591
R545 avss.n146 avss.n145 53.0711
R546 avss.n47 avss.n43 52.8748
R547 avss.n323 avss.t135 51.2742
R548 avss.n155 avss.t41 50.6958
R549 avss.n139 avss.t119 43.7033
R550 avss.n299 avss.t39 40.2071
R551 avss.n345 avss.n344 37.0713
R552 avss.n181 avss.t24 36.7109
R553 avss.n38 avss.t78 34.5898
R554 avss.t98 avss.t132 34.0887
R555 avss.t16 avss.t142 34.0887
R556 avss.n145 avss.n51 33.6939
R557 avss.n296 avss.n51 33.6822
R558 avss.n222 avss.t128 33.2146
R559 avss.n289 avss.t149 31.4665
R560 avss.n312 avss.n311 31.4345
R561 avss.n312 avss.n42 31.1137
R562 avss.t162 avss.t29 30.5925
R563 avss.n219 avss.t51 29.7184
R564 avss.t12 avss.t66 27.0962
R565 avss.n177 avss.t144 26.2222
R566 avss.n127 avss.t43 24.4741
R567 avss.t6 avss.t83 23.6
R568 avss.n293 avss.n51 23.2228
R569 avss.n158 avss.n61 22.7741
R570 avss.n161 avss.n159 22.7741
R571 avss.n161 avss.n160 22.7741
R572 avss.n257 avss.n76 22.7741
R573 avss.n257 avss.n256 22.7741
R574 avss.n255 avss.n254 22.7741
R575 avss.n254 avss.n79 22.7741
R576 avss.n188 avss.n186 22.7741
R577 avss.n188 avss.n187 22.7741
R578 avss.n239 avss.n100 22.7741
R579 avss.n239 avss.n238 22.7741
R580 avss.n237 avss.n236 22.7741
R581 avss.n236 avss.n103 22.7741
R582 avss.n213 avss.n211 22.7741
R583 avss.n213 avss.n212 22.7741
R584 avss.n147 avss.n146 22.7741
R585 avss.n149 avss.n148 22.7741
R586 avss.n150 avss.n149 22.7741
R587 avss.n164 avss.n131 22.7741
R588 avss.n165 avss.n164 22.7741
R589 avss.n167 avss.n166 22.7741
R590 avss.n168 avss.n167 22.7741
R591 avss.n170 avss.n169 22.7741
R592 avss.n191 avss.n119 22.7741
R593 avss.n192 avss.n191 22.7741
R594 avss.n194 avss.n193 22.7741
R595 avss.n195 avss.n194 22.7741
R596 avss.n197 avss.n196 22.7741
R597 avss.n198 avss.n197 22.7741
R598 avss.n207 avss.n199 22.7741
R599 avss.n207 avss.n206 22.7741
R600 avss.n205 avss.n204 22.7741
R601 avss.n328 avss.n7 22.6318
R602 avss.n330 avss.n24 22.6318
R603 avss.n330 avss.n329 22.6318
R604 avss.n26 avss.n8 22.3524
R605 avss.n334 avss.n333 22.3524
R606 avss.n225 avss.n13 22.0798
R607 avss.n233 avss.n108 22.0798
R608 avss.n243 avss.n242 22.0798
R609 avss.n184 avss.n90 22.0798
R610 avss.n251 avss.n84 22.0798
R611 avss.n261 avss.n260 22.0798
R612 avss.n142 avss.n66 22.0798
R613 avss.n155 avss.n154 21.8519
R614 avss.n27 avss.t122 20.9779
R615 avss.n286 avss.n61 20.9565
R616 avss.n313 avss.n312 20.857
R617 avss.n295 avss.n294 20.8255
R618 avss.n286 avss.n285 20.3176
R619 avss.n294 avss.n293 20.3176
R620 avss.t4 avss.t59 20.1038
R621 avss.n324 avss.t115 20.1038
R622 avss.n307 avss.n306 20.0728
R623 avss.n306 avss.n304 19.868
R624 avss.n172 avss.n170 19.2458
R625 avss.t48 avss.n153 19.2297
R626 avss.n270 avss.n269 18.2614
R627 avss.n36 avss.n31 18.2614
R628 avss.n322 avss.n321 18.2614
R629 avss.n349 avss.n348 18.2614
R630 avss.n305 avss.n41 18.1811
R631 avss.n115 avss.t166 17.4816
R632 avss.n344 avss.n8 16.8713
R633 avss.t10 avss.t147 16.6076
R634 avss.n116 avss.t61 13.9854
R635 avss.n159 avss.n158 13.8999
R636 avss.n160 avss.n76 13.8999
R637 avss.n256 avss.n255 13.8999
R638 avss.n186 avss.n79 13.8999
R639 avss.n187 avss.n100 13.8999
R640 avss.n238 avss.n237 13.8999
R641 avss.n211 avss.n103 13.8999
R642 avss.n150 avss.n131 13.8999
R643 avss.n166 avss.n165 13.8999
R644 avss.n169 avss.n168 13.8999
R645 avss.n173 avss.n119 13.8999
R646 avss.n193 avss.n192 13.8999
R647 avss.n196 avss.n195 13.8999
R648 avss.n199 avss.n198 13.8999
R649 avss.n206 avss.n205 13.8999
R650 avss.n212 avss.n24 13.8885
R651 avss.n329 avss.n328 13.8772
R652 avss.n333 avss.n20 13.8524
R653 avss.n201 avss.n26 13.8326
R654 avss.n335 avss.n334 13.8108
R655 avss.n226 avss.n225 13.789
R656 avss.n113 avss.n108 13.789
R657 avss.n244 avss.n243 13.789
R658 avss.n184 avss.n86 13.789
R659 avss.n125 avss.n84 13.789
R660 avss.n262 avss.n261 13.789
R661 avss.n142 avss.n63 13.789
R662 avss.n336 avss.n13 13.6834
R663 avss.n233 avss.n232 13.6834
R664 avss.n242 avss.n96 13.6834
R665 avss.n245 avss.n90 13.6834
R666 avss.n251 avss.n250 13.6834
R667 avss.n260 avss.n72 13.6834
R668 avss.n263 avss.n66 13.6834
R669 avss.n285 avss.n284 13.6834
R670 avss.n60 avss.n53 13.0308
R671 avss.n171 avss.n89 11.2624
R672 avss.n171 avss.n65 10.8741
R673 avss.n325 avss.t114 10.4892
R674 avss.t18 avss.t63 9.61512
R675 avss.n268 avss.n267 8.67882
R676 avss.n201 avss.n20 8.5005
R677 avss.n336 avss.n335 8.39684
R678 avss.n232 avss.n226 8.39684
R679 avss.n113 avss.n96 8.39684
R680 avss.n245 avss.n244 8.39684
R681 avss.n250 avss.n86 8.39684
R682 avss.n125 avss.n72 8.39684
R683 avss.n263 avss.n262 8.39684
R684 avss.n284 avss.n63 8.39684
R685 avss.n341 avss.n11 7.576
R686 avss.n298 avss.t80 6.99295
R687 avss.n128 avss.t54 6.99295
R688 avss.n287 avss.n60 6.57174
R689 avss.n64 avss.n60 5.75386
R690 avss.n344 avss.n343 5.7505
R691 avss.n47 avss.n46 5.7505
R692 avss.n303 avss.n34 5.7505
R693 avss.n320 avss.n29 5.06074
R694 avss.n37 avss.n29 5.06074
R695 avss.n30 avss.n28 5.06074
R696 avss.n37 avss.n28 5.06074
R697 avss.n4 avss.n2 5.06074
R698 avss.n154 avss.n4 5.06074
R699 avss.n267 avss.n3 5.06074
R700 avss.n154 avss.n3 5.06074
R701 avss.n306 avss.n305 5.03754
R702 avss.n278 avss.n277 4.24397
R703 avss.n271 avss.n270 4.08577
R704 avss.n275 avss.n273 4.02904
R705 avss.n278 avss.n276 4.02846
R706 avss.n350 avss.n349 3.86414
R707 avss.n343 avss.n342 3.7505
R708 avss.n173 avss.n172 3.5288
R709 avss.n337 avss.n336 2.8755
R710 avss.n232 avss.n231 2.8755
R711 avss.n227 avss.n96 2.8755
R712 avss.n246 avss.n245 2.8755
R713 avss.n250 avss.n249 2.8755
R714 avss.n87 avss.n72 2.8755
R715 avss.n264 avss.n263 2.8755
R716 avss.n284 avss.n283 2.8755
R717 avss.n20 avss.n19 2.8755
R718 avss.n305 avss.n32 2.55606
R719 avss.n10 avss 2.41717
R720 avss.n274 avss.n273 2.28395
R721 avss.n282 avss.n64 1.92646
R722 avss.n19 avss.n9 1.8755
R723 avss.n228 avss.n227 1.8755
R724 avss.n231 avss.n230 1.8755
R725 avss.n338 avss.n337 1.8755
R726 avss.n88 avss.n87 1.8755
R727 avss.n249 avss.n248 1.8755
R728 avss.n247 avss.n246 1.8755
R729 avss.n283 avss.n282 1.8755
R730 avss.n265 avss.n264 1.8755
R731 avss.n307 avss.n47 1.84387
R732 avss.n229 avss.n1 1.57742
R733 avss.n268 avss.n266 1.57742
R734 avss.n351 avss.n350 1.35235
R735 avss.n272 avss.n271 1.35235
R736 avss.n304 avss.n303 1.22942
R737 avss.n319 avss.n318 1.1505
R738 avss.n340 avss.n339 0.465313
R739 avss.n281 avss.n272 0.413757
R740 avss.n172 avss.n171 0.392043
R741 avss.n287 avss.n286 0.381766
R742 avss.n340 avss.n0 0.352634
R743 avss.n342 avss.n9 0.282818
R744 avss.n248 avss.n88 0.267454
R745 avss.n248 avss.n247 0.267454
R746 avss.n247 avss.n89 0.236725
R747 avss.n294 avss.n53 0.216817
R748 avss.n279 avss.n278 0.215807
R749 avss.n280 avss.n12 0.189131
R750 avss.n313 avss.n41 0.157907
R751 avss.n341 avss.n340 0.148664
R752 avss avss.n351 0.123411
R753 avss.n88 avss.n65 0.121013
R754 avss.n12 avss.n0 0.110668
R755 avss.n11 avss.n10 0.0793127
R756 avss.n281 avss.n280 0.0674007
R757 avss.n46 avss.n32 0.056753
R758 avss.n230 avss.n228 0.0514608
R759 avss.n280 avss.n279 0.0489848
R760 avss.n266 avss.n265 0.0484362
R761 avss.n339 avss.n338 0.0447699
R762 avss.n10 avss 0.0387586
R763 avss.n317 avss.n34 0.037012
R764 avss.t110 avss.n274 0.0366713
R765 avss.n339 avss.n9 0.0355497
R766 avss.n338 avss.n12 0.032213
R767 avss.n265 avss.n65 0.0284551
R768 avss.t31 avss.n275 0.025875
R769 avss.t36 avss.n276 0.025875
R770 avss.n277 avss.t44 0.025875
R771 avss.n275 avss.t110 0.0217625
R772 avss.n276 avss.t31 0.0217625
R773 avss.n277 avss.t36 0.0217625
R774 avss.n230 avss.n229 0.0196561
R775 avss.n34 avss.n33 0.0190181
R776 avss.n318 avss.n32 0.0186687
R777 avss.n342 avss.n341 0.0125033
R778 avss.n274 avss.t164 0.0119119
R779 avss.n33 avss.n11 0.00783735
R780 avss.n228 avss.n89 0.00636599
R781 avss.n272 avss 0.00391775
R782 avss.n282 avss.n281 0.003433
R783 avss.n279 avss.n273 0.000702166
R784 avss.n318 avss.n317 0.000674699
R785 avss.n351 avss.n0 0.000623404
R786 avss.n229 avss.n12 0.000591656
R787 avss.n281 avss.n266 0.000591656
R788 ena.n5 ena.t2 546.938
R789 ena.n5 ena.t3 530.298
R790 ena.n1 ena.t5 446.656
R791 ena.n0 ena.t6 442.243
R792 ena.n3 ena.t4 310.555
R793 ena.n2 ena.t1 181.511
R794 ena.n2 ena.t0 177.388
R795 ena.n5 ena.n4 15.0005
R796 ena.n4 ena.n3 2.36247
R797 ena.n4 ena.n1 1.99822
R798 ena.n3 ena.n2 1.39855
R799 ena.n1 ena.n0 1.23837
R800 ena.n0 ena 0.427444
R801 ena ena.n5 0.072275
R802 avdd.n245 avdd.n244 46118
R803 avdd.n244 avdd.n230 46118
R804 avdd.n246 avdd.n245 32152.6
R805 avdd.n298 avdd.n230 32148.4
R806 avdd.n243 avdd.n228 19114.5
R807 avdd.n243 avdd.n240 19114.5
R808 avdd.n247 avdd.n240 13442.8
R809 avdd.n299 avdd.n228 13441.1
R810 avdd.n298 avdd.n297 11487.6
R811 avdd.n246 avdd.n231 11466.6
R812 avdd.n297 avdd.n296 8703.73
R813 avdd.n299 avdd.n229 5050.22
R814 avdd.n248 avdd.n247 5041.7
R815 avdd.n296 avdd.n231 5039.44
R816 avdd.n248 avdd.n232 4168.22
R817 avdd.n232 avdd.n229 4161.41
R818 avdd.n242 avdd.n241 1663.09
R819 avdd.n226 avdd.n0 1347.44
R820 avdd.n241 avdd.n239 1260.78
R821 avdd.n301 avdd.n226 1006.53
R822 avdd.n167 avdd.t22 942.102
R823 avdd.n167 avdd.t15 942.087
R824 avdd.n5 avdd.t3 942.087
R825 avdd.n94 avdd.t5 942.087
R826 avdd.n106 avdd.t9 942.087
R827 avdd.n165 avdd.t7 942.087
R828 avdd.n221 avdd.t11 942.087
R829 avdd.n4 avdd.t1 942.087
R830 avdd.n206 avdd.t13 942.087
R831 avdd.n253 avdd.t17 941.889
R832 avdd.n290 avdd.t20 941.876
R833 avdd.n154 avdd.n144 929.793
R834 avdd.n154 avdd.n145 929.793
R835 avdd.n144 avdd.n143 929.793
R836 avdd.n145 avdd.n143 929.793
R837 avdd.n172 avdd.n120 929.793
R838 avdd.n172 avdd.n121 929.793
R839 avdd.n171 avdd.n121 929.793
R840 avdd.n171 avdd.n120 929.793
R841 avdd.n177 avdd.n114 929.793
R842 avdd.n177 avdd.n115 929.793
R843 avdd.n115 avdd.n113 929.793
R844 avdd.n114 avdd.n113 929.793
R845 avdd.n196 avdd.n87 929.793
R846 avdd.n185 avdd.n87 929.793
R847 avdd.n185 avdd.n88 929.793
R848 avdd.n196 avdd.n88 929.793
R849 avdd.n201 avdd.n83 929.793
R850 avdd.n199 avdd.n83 929.793
R851 avdd.n200 avdd.n199 929.793
R852 avdd.n201 avdd.n200 929.793
R853 avdd.n211 avdd.n21 929.793
R854 avdd.n211 avdd.n22 929.793
R855 avdd.n210 avdd.n22 929.793
R856 avdd.n210 avdd.n21 929.793
R857 avdd.n216 avdd.n17 929.793
R858 avdd.n216 avdd.n18 929.793
R859 avdd.n18 avdd.n11 929.793
R860 avdd.n17 avdd.n11 929.793
R861 avdd.n141 avdd.n139 929.793
R862 avdd.n155 avdd.n139 929.793
R863 avdd.n155 avdd.n138 929.793
R864 avdd.n141 avdd.n138 929.793
R865 avdd.n128 avdd.n123 929.793
R866 avdd.n128 avdd.n124 929.793
R867 avdd.n134 avdd.n124 929.793
R868 avdd.n134 avdd.n123 929.793
R869 avdd.n110 avdd.n109 929.793
R870 avdd.n178 avdd.n110 929.793
R871 avdd.n179 avdd.n178 929.793
R872 avdd.n179 avdd.n109 929.793
R873 avdd.n187 avdd.n99 929.793
R874 avdd.n188 avdd.n187 929.793
R875 avdd.n188 avdd.n86 929.793
R876 avdd.n99 avdd.n86 929.793
R877 avdd.n85 avdd.n81 929.793
R878 avdd.n85 avdd.n82 929.793
R879 avdd.n203 avdd.n82 929.793
R880 avdd.n203 avdd.n81 929.793
R881 avdd.n28 avdd.n24 929.793
R882 avdd.n28 avdd.n25 929.793
R883 avdd.n32 avdd.n25 929.793
R884 avdd.n32 avdd.n24 929.793
R885 avdd.n217 avdd.n13 929.793
R886 avdd.n15 avdd.n13 929.793
R887 avdd.n15 avdd.n12 929.793
R888 avdd.n217 avdd.n12 929.793
R889 avdd.n56 avdd.n49 929.793
R890 avdd.n53 avdd.n49 929.793
R891 avdd.n56 avdd.n48 929.793
R892 avdd.n70 avdd.n43 929.793
R893 avdd.n70 avdd.n44 929.793
R894 avdd.n43 avdd.n42 929.793
R895 avdd.n44 avdd.n42 929.793
R896 avdd.n40 avdd.n37 929.793
R897 avdd.n40 avdd.n38 929.793
R898 avdd.n71 avdd.n38 929.793
R899 avdd.n71 avdd.n37 929.793
R900 avdd.n266 avdd.n264 929.793
R901 avdd.n275 avdd.n264 929.793
R902 avdd.n275 avdd.n269 929.793
R903 avdd.n269 avdd.n266 929.793
R904 avdd.n285 avdd.n256 929.793
R905 avdd.n286 avdd.n256 929.793
R906 avdd.n285 avdd.n257 929.793
R907 avdd.n286 avdd.n257 929.793
R908 avdd.n272 avdd.n234 929.793
R909 avdd.n272 avdd.n235 929.793
R910 avdd.n294 avdd.n235 929.793
R911 avdd.n294 avdd.n234 929.793
R912 avdd.n277 avdd.n259 929.793
R913 avdd.n281 avdd.n259 929.793
R914 avdd.n277 avdd.n260 929.793
R915 avdd.n281 avdd.n260 929.793
R916 avdd.n249 avdd.n239 449.079
R917 avdd.n55 avdd.n39 442.036
R918 avdd.n300 avdd.n227 405.76
R919 avdd.n250 avdd.n249 305.716
R920 avdd.n296 avdd.n295 239.046
R921 avdd.n251 avdd.n238 238.297
R922 avdd.t23 avdd.n55 212.059
R923 avdd.t2 avdd.n39 212.059
R924 avdd.t2 avdd.n41 212.059
R925 avdd.t0 avdd.n14 212.059
R926 avdd.t0 avdd.n16 212.059
R927 avdd.t10 avdd.n23 212.059
R928 avdd.t10 avdd.n26 212.059
R929 avdd.n202 avdd.t12 212.059
R930 avdd.n198 avdd.t12 212.059
R931 avdd.n197 avdd.t4 212.059
R932 avdd.n186 avdd.t4 212.059
R933 avdd.t8 avdd.n101 212.059
R934 avdd.t8 avdd.n112 212.059
R935 avdd.t6 avdd.n122 212.059
R936 avdd.t6 avdd.n125 212.059
R937 avdd.t14 avdd.n140 212.059
R938 avdd.t14 avdd.n142 212.059
R939 avdd.n54 avdd.n48 196.584
R940 avdd.n41 avdd.n14 189.16
R941 avdd.n23 avdd.n16 189.16
R942 avdd.n202 avdd.n26 189.16
R943 avdd.n198 avdd.n197 189.16
R944 avdd.n186 avdd.n101 189.16
R945 avdd.n122 avdd.n112 189.16
R946 avdd.n140 avdd.n125 189.16
R947 avdd.t18 avdd.n258 183.154
R948 avdd.t18 avdd.n261 183.154
R949 avdd.t16 avdd.n233 177.994
R950 avdd.n273 avdd.t21 177.994
R951 avdd.n274 avdd.n258 158.218
R952 avdd.n147 avdd.n137 151.554
R953 avdd.n152 avdd.n147 149.745
R954 avdd.n135 avdd.n126 122.114
R955 avdd.n181 avdd.n180 122.114
R956 avdd.n97 avdd.n95 122.114
R957 avdd.n33 avdd.n7 122.114
R958 avdd.n34 avdd.n10 122.114
R959 avdd.n62 avdd.n61 122.114
R960 avdd.n136 avdd.n131 122.114
R961 avdd.n205 avdd.n204 122.114
R962 avdd.n207 avdd.n30 119.614
R963 avdd.n164 avdd.n118 119.614
R964 avdd.n182 avdd.n105 119.614
R965 avdd.n195 avdd.n194 119.614
R966 avdd.n220 avdd.n6 119.614
R967 avdd.n65 avdd.n64 119.614
R968 avdd.n60 avdd.n59 119.614
R969 avdd.n168 avdd.n130 119.614
R970 avdd.n169 avdd.n129 113.501
R971 avdd.n163 avdd.n162 113.501
R972 avdd.n183 avdd.n100 113.501
R973 avdd.n193 avdd.n192 113.501
R974 avdd.n208 avdd.n29 113.501
R975 avdd.n219 avdd.n9 113.501
R976 avdd.n58 avdd.n46 113.501
R977 avdd.n66 avdd.n35 113.501
R978 avdd.n158 avdd.n129 113.001
R979 avdd.n160 avdd.n135 113.001
R980 avdd.n162 avdd.n161 113.001
R981 avdd.n180 avdd.n108 113.001
R982 avdd.n100 avdd.n98 113.001
R983 avdd.n190 avdd.n97 113.001
R984 avdd.n192 avdd.n191 113.001
R985 avdd.n79 avdd.n29 113.001
R986 avdd.n77 avdd.n33 113.001
R987 avdd.n74 avdd.n34 113.001
R988 avdd.n76 avdd.n9 113.001
R989 avdd.n51 avdd.n46 113.001
R990 avdd.n73 avdd.n35 113.001
R991 avdd.n61 avdd.n36 113.001
R992 avdd.n157 avdd.n136 113.001
R993 avdd.n204 avdd.n80 113.001
R994 avdd.n169 avdd.n127 111.501
R995 avdd.n163 avdd.n117 111.501
R996 avdd.n184 avdd.n183 111.501
R997 avdd.n193 avdd.n84 111.501
R998 avdd.n208 avdd.n27 111.501
R999 avdd.n219 avdd.n8 111.501
R1000 avdd.n67 avdd.n66 111.501
R1001 avdd.n89 avdd.n30 110.001
R1002 avdd.n127 avdd.n119 110.001
R1003 avdd.n174 avdd.n118 110.001
R1004 avdd.n175 avdd.n117 110.001
R1005 avdd.n116 avdd.n105 110.001
R1006 avdd.n184 avdd.n103 110.001
R1007 avdd.n195 avdd.n93 110.001
R1008 avdd.n92 avdd.n84 110.001
R1009 avdd.n27 avdd.n20 110.001
R1010 avdd.n213 avdd.n6 110.001
R1011 avdd.n64 avdd.n19 110.001
R1012 avdd.n214 avdd.n8 110.001
R1013 avdd.n68 avdd.n67 110.001
R1014 avdd.n59 avdd.n45 110.001
R1015 avdd.n146 avdd.n130 110.001
R1016 avdd.n47 avdd.n45 85.6283
R1017 avdd.n57 avdd.n56 70.0005
R1018 avdd.n56 avdd.t23 70.0005
R1019 avdd.n218 avdd.n217 70.0005
R1020 avdd.n217 avdd.t0 70.0005
R1021 avdd.n209 avdd.n24 70.0005
R1022 avdd.t10 avdd.n24 70.0005
R1023 avdd.n81 avdd.n31 70.0005
R1024 avdd.t12 avdd.n81 70.0005
R1025 avdd.n104 avdd.n99 70.0005
R1026 avdd.n99 avdd.t4 70.0005
R1027 avdd.n109 avdd.n107 70.0005
R1028 avdd.t8 avdd.n109 70.0005
R1029 avdd.n170 avdd.n123 70.0005
R1030 avdd.t6 avdd.n123 70.0005
R1031 avdd.n149 avdd.n141 70.0005
R1032 avdd.t14 avdd.n141 70.0005
R1033 avdd.n218 avdd.n11 70.0005
R1034 avdd.t0 avdd.n11 70.0005
R1035 avdd.n210 avdd.n209 70.0005
R1036 avdd.t10 avdd.n210 70.0005
R1037 avdd.n200 avdd.n31 70.0005
R1038 avdd.n200 avdd.t12 70.0005
R1039 avdd.n104 avdd.n88 70.0005
R1040 avdd.n88 avdd.t4 70.0005
R1041 avdd.n113 avdd.n107 70.0005
R1042 avdd.t8 avdd.n113 70.0005
R1043 avdd.n171 avdd.n170 70.0005
R1044 avdd.t6 avdd.n171 70.0005
R1045 avdd.n149 avdd.n143 70.0005
R1046 avdd.t14 avdd.n143 70.0005
R1047 avdd.n63 avdd.n42 70.0005
R1048 avdd.t2 avdd.n42 70.0005
R1049 avdd.n63 avdd.n40 70.0005
R1050 avdd.t2 avdd.n40 70.0005
R1051 avdd.n70 avdd.n69 70.0005
R1052 avdd.t2 avdd.n70 70.0005
R1053 avdd.n216 avdd.n215 70.0005
R1054 avdd.t0 avdd.n216 70.0005
R1055 avdd.n212 avdd.n211 70.0005
R1056 avdd.n211 avdd.t10 70.0005
R1057 avdd.n91 avdd.n83 70.0005
R1058 avdd.n83 avdd.t12 70.0005
R1059 avdd.n102 avdd.n87 70.0005
R1060 avdd.n87 avdd.t4 70.0005
R1061 avdd.n177 avdd.n176 70.0005
R1062 avdd.t8 avdd.n177 70.0005
R1063 avdd.n173 avdd.n172 70.0005
R1064 avdd.n172 avdd.t6 70.0005
R1065 avdd.n154 avdd.n153 70.0005
R1066 avdd.t14 avdd.n154 70.0005
R1067 avdd.n53 avdd.n52 70.0005
R1068 avdd.n72 avdd.n71 70.0005
R1069 avdd.n71 avdd.t2 70.0005
R1070 avdd.n75 avdd.n15 70.0005
R1071 avdd.t0 avdd.n15 70.0005
R1072 avdd.n78 avdd.n25 70.0005
R1073 avdd.t10 avdd.n25 70.0005
R1074 avdd.n96 avdd.n82 70.0005
R1075 avdd.t12 avdd.n82 70.0005
R1076 avdd.n189 avdd.n188 70.0005
R1077 avdd.n188 avdd.t4 70.0005
R1078 avdd.n178 avdd.n111 70.0005
R1079 avdd.n178 avdd.t8 70.0005
R1080 avdd.n159 avdd.n124 70.0005
R1081 avdd.t6 avdd.n124 70.0005
R1082 avdd.n156 avdd.n155 70.0005
R1083 avdd.n155 avdd.t14 70.0005
R1084 avdd.n267 avdd.n234 70.0005
R1085 avdd.t16 avdd.n234 70.0005
R1086 avdd.n237 avdd.n235 70.0005
R1087 avdd.t16 avdd.n235 70.0005
R1088 avdd.n287 avdd.n286 70.0005
R1089 avdd.n286 avdd.t18 70.0005
R1090 avdd.n269 avdd.n268 70.0005
R1091 avdd.t21 avdd.n269 70.0005
R1092 avdd.n280 avdd.n259 70.0005
R1093 avdd.t18 avdd.n259 70.0005
R1094 avdd.n264 avdd.n263 70.0005
R1095 avdd.t21 avdd.n264 70.0005
R1096 avdd.n285 avdd.n284 70.0005
R1097 avdd.t18 avdd.n285 70.0005
R1098 avdd.n284 avdd.n260 70.0005
R1099 avdd.t18 avdd.n260 70.0005
R1100 avdd.n265 avdd.n263 67.907
R1101 avdd.n282 avdd.n280 66.9661
R1102 avdd.n242 avdd.n0 66.0812
R1103 avdd.n52 avdd.n50 59.6701
R1104 avdd.n50 avdd.n48 56.0005
R1105 avdd.n49 avdd.n46 56.0005
R1106 avdd.n55 avdd.n49 56.0005
R1107 avdd.n34 avdd.n12 56.0005
R1108 avdd.n14 avdd.n12 56.0005
R1109 avdd.n13 avdd.n9 56.0005
R1110 avdd.n16 avdd.n13 56.0005
R1111 avdd.n33 avdd.n32 56.0005
R1112 avdd.n32 avdd.n23 56.0005
R1113 avdd.n29 avdd.n28 56.0005
R1114 avdd.n28 avdd.n26 56.0005
R1115 avdd.n192 avdd.n85 56.0005
R1116 avdd.n198 avdd.n85 56.0005
R1117 avdd.n97 avdd.n86 56.0005
R1118 avdd.n197 avdd.n86 56.0005
R1119 avdd.n187 avdd.n100 56.0005
R1120 avdd.n187 avdd.n186 56.0005
R1121 avdd.n180 avdd.n179 56.0005
R1122 avdd.n179 avdd.n101 56.0005
R1123 avdd.n162 avdd.n110 56.0005
R1124 avdd.n112 avdd.n110 56.0005
R1125 avdd.n135 avdd.n134 56.0005
R1126 avdd.n134 avdd.n122 56.0005
R1127 avdd.n129 avdd.n128 56.0005
R1128 avdd.n128 avdd.n125 56.0005
R1129 avdd.n148 avdd.n139 56.0005
R1130 avdd.n142 avdd.n139 56.0005
R1131 avdd.n64 avdd.n17 56.0005
R1132 avdd.n17 avdd.n14 56.0005
R1133 avdd.n18 avdd.n8 56.0005
R1134 avdd.n18 avdd.n16 56.0005
R1135 avdd.n21 avdd.n6 56.0005
R1136 avdd.n23 avdd.n21 56.0005
R1137 avdd.n27 avdd.n22 56.0005
R1138 avdd.n26 avdd.n22 56.0005
R1139 avdd.n201 avdd.n30 56.0005
R1140 avdd.n202 avdd.n201 56.0005
R1141 avdd.n199 avdd.n84 56.0005
R1142 avdd.n199 avdd.n198 56.0005
R1143 avdd.n196 avdd.n195 56.0005
R1144 avdd.n197 avdd.n196 56.0005
R1145 avdd.n185 avdd.n184 56.0005
R1146 avdd.n186 avdd.n185 56.0005
R1147 avdd.n114 avdd.n105 56.0005
R1148 avdd.n114 avdd.n101 56.0005
R1149 avdd.n117 avdd.n115 56.0005
R1150 avdd.n115 avdd.n112 56.0005
R1151 avdd.n120 avdd.n118 56.0005
R1152 avdd.n122 avdd.n120 56.0005
R1153 avdd.n127 avdd.n121 56.0005
R1154 avdd.n125 avdd.n121 56.0005
R1155 avdd.n151 avdd.n145 56.0005
R1156 avdd.n145 avdd.n142 56.0005
R1157 avdd.n67 avdd.n44 56.0005
R1158 avdd.n44 avdd.n41 56.0005
R1159 avdd.n38 avdd.n35 56.0005
R1160 avdd.n41 avdd.n38 56.0005
R1161 avdd.n61 avdd.n37 56.0005
R1162 avdd.n39 avdd.n37 56.0005
R1163 avdd.n59 avdd.n43 56.0005
R1164 avdd.n43 avdd.n39 56.0005
R1165 avdd.n144 avdd.n130 56.0005
R1166 avdd.n144 avdd.n140 56.0005
R1167 avdd.n138 avdd.n136 56.0005
R1168 avdd.n140 avdd.n138 56.0005
R1169 avdd.n204 avdd.n203 56.0005
R1170 avdd.n203 avdd.n202 56.0005
R1171 avdd.n294 avdd.n293 56.0005
R1172 avdd.n295 avdd.n294 56.0005
R1173 avdd.n266 avdd.n265 56.0005
R1174 avdd.n266 avdd.n233 56.0005
R1175 avdd.n282 avdd.n281 56.0005
R1176 avdd.n281 avdd.n261 56.0005
R1177 avdd.n276 avdd.n275 56.0005
R1178 avdd.n275 avdd.n274 56.0005
R1179 avdd.n278 avdd.n277 56.0005
R1180 avdd.n277 avdd.n258 56.0005
R1181 avdd.n272 avdd.n271 56.0005
R1182 avdd.n273 avdd.n272 56.0005
R1183 avdd.n271 avdd.n256 56.0005
R1184 avdd.n258 avdd.n256 56.0005
R1185 avdd.n257 avdd.n254 56.0005
R1186 avdd.n261 avdd.n257 56.0005
R1187 avdd.n156 avdd.n137 52.9895
R1188 avdd.n50 avdd.n47 52.5666
R1189 avdd.n153 avdd.n152 52.1466
R1190 avdd.n54 avdd.n53 51.3363
R1191 avdd.n296 avdd.n232 51.0335
R1192 avdd.n51 avdd.n36 47.4722
R1193 avdd.n288 avdd.n287 35.3541
R1194 avdd.n292 avdd.n237 34.4183
R1195 avdd.n238 avdd.n227 33.4758
R1196 avdd.n60 avdd.n58 32.0925
R1197 avdd.n150 avdd.n148 31.8931
R1198 avdd.n151 avdd.n150 31.3311
R1199 avdd.n280 avdd.n279 30.8524
R1200 avdd.n279 avdd.n263 30.8524
R1201 avdd.n293 avdd.n236 30.7069
R1202 avdd.n293 avdd.n292 30.6275
R1203 avdd.n283 avdd.n282 30.6275
R1204 avdd.n283 avdd.n254 30.6275
R1205 avdd.n265 avdd.n236 30.1489
R1206 avdd.n288 avdd.n254 29.1434
R1207 avdd.n287 avdd.n255 26.8715
R1208 avdd.n255 avdd.n237 26.8715
R1209 avdd.n271 avdd.n262 25.3487
R1210 avdd.n69 avdd.n45 22.7741
R1211 avdd.n69 avdd.n68 22.7741
R1212 avdd.n215 avdd.n19 22.7741
R1213 avdd.n215 avdd.n214 22.7741
R1214 avdd.n213 avdd.n212 22.7741
R1215 avdd.n212 avdd.n20 22.7741
R1216 avdd.n92 avdd.n91 22.7741
R1217 avdd.n102 avdd.n93 22.7741
R1218 avdd.n103 avdd.n102 22.7741
R1219 avdd.n176 avdd.n116 22.7741
R1220 avdd.n176 avdd.n175 22.7741
R1221 avdd.n174 avdd.n173 22.7741
R1222 avdd.n173 avdd.n119 22.7741
R1223 avdd.n153 avdd.n146 22.7741
R1224 avdd.n52 avdd.n51 22.7741
R1225 avdd.n72 avdd.n36 22.7741
R1226 avdd.n73 avdd.n72 22.7741
R1227 avdd.n75 avdd.n74 22.7741
R1228 avdd.n76 avdd.n75 22.7741
R1229 avdd.n78 avdd.n77 22.7741
R1230 avdd.n79 avdd.n78 22.7741
R1231 avdd.n96 avdd.n80 22.7741
R1232 avdd.n191 avdd.n96 22.7741
R1233 avdd.n190 avdd.n189 22.7741
R1234 avdd.n189 avdd.n98 22.7741
R1235 avdd.n111 avdd.n108 22.7741
R1236 avdd.n161 avdd.n111 22.7741
R1237 avdd.n160 avdd.n159 22.7741
R1238 avdd.n159 avdd.n158 22.7741
R1239 avdd.n157 avdd.n156 22.7741
R1240 avdd.n279 avdd.n278 21.6014
R1241 avdd.n68 avdd.n19 20.315
R1242 avdd.n214 avdd.n213 20.315
R1243 avdd.n89 avdd.n20 20.315
R1244 avdd.n93 avdd.n92 20.315
R1245 avdd.n116 avdd.n103 20.315
R1246 avdd.n175 avdd.n174 20.315
R1247 avdd.n146 avdd.n119 20.315
R1248 avdd.n74 avdd.n73 20.315
R1249 avdd.n77 avdd.n76 20.315
R1250 avdd.n80 avdd.n79 20.315
R1251 avdd.n191 avdd.n190 20.315
R1252 avdd.n108 avdd.n98 20.315
R1253 avdd.n161 avdd.n160 20.315
R1254 avdd.n158 avdd.n157 20.315
R1255 avdd.n267 avdd.n236 20.1781
R1256 avdd.n284 avdd.n283 19.7551
R1257 avdd.n150 avdd.n149 19.1628
R1258 avdd.n276 avdd.n262 17.6244
R1259 avdd.n170 avdd.n169 15.8821
R1260 avdd.n163 avdd.n107 15.8821
R1261 avdd.n183 avdd.n104 15.8821
R1262 avdd.n193 avdd.n31 15.8821
R1263 avdd.n209 avdd.n208 15.8821
R1264 avdd.n219 avdd.n218 15.8821
R1265 avdd.n66 avdd.n63 15.8821
R1266 avdd.n58 avdd.n57 15.8446
R1267 avdd.n284 avdd.n262 15.4264
R1268 avdd.n268 avdd.n262 15.094
R1269 avdd.t23 avdd.n54 14.8009
R1270 avdd.n90 avdd.n89 14.4345
R1271 avdd.n169 avdd.n168 12.9863
R1272 avdd.n164 avdd.n163 12.9863
R1273 avdd.n183 avdd.n182 12.9863
R1274 avdd.n194 avdd.n193 12.9863
R1275 avdd.n208 avdd.n207 12.9863
R1276 avdd.n220 avdd.n219 12.9863
R1277 avdd.n66 avdd.n65 12.9863
R1278 avdd.n271 avdd.n270 11.688
R1279 avdd.n148 avdd.n137 10.9592
R1280 avdd.n152 avdd.n151 10.8187
R1281 avdd.n270 avdd.n255 10.0943
R1282 avdd.n249 avdd.n248 9.33383
R1283 avdd.n248 avdd.n231 9.33383
R1284 avdd.n229 avdd.n227 9.33383
R1285 avdd.n297 avdd.n229 9.33383
R1286 avdd.n91 avdd.n90 8.34012
R1287 avdd.n289 avdd.n288 7.67637
R1288 avdd.n292 avdd.n291 7.66717
R1289 avdd.n250 avdd.n232 7.17999
R1290 avdd.n295 avdd.n233 5.15974
R1291 avdd.t21 avdd.t16 5.15974
R1292 avdd.n274 avdd.n273 5.15974
R1293 avdd.n247 avdd.n239 5.09141
R1294 avdd.n247 avdd.n246 5.09141
R1295 avdd.n300 avdd.n299 5.09141
R1296 avdd.n299 avdd.n298 5.09141
R1297 avdd.n150 avdd.n147 4.47418
R1298 avdd.n251 avdd.n250 3.42332
R1299 avdd.n57 avdd.n47 3.34111
R1300 avdd.n270 avdd.n253 2.3005
R1301 avdd.n165 avdd.n164 1.91717
R1302 avdd.n182 avdd.n106 1.91717
R1303 avdd.n194 avdd.n94 1.91717
R1304 avdd.n221 avdd.n220 1.91717
R1305 avdd.n65 avdd.n4 1.91717
R1306 avdd.n60 avdd.n5 1.91717
R1307 avdd.n168 avdd.n167 1.91717
R1308 avdd.n207 avdd.n206 1.91717
R1309 avdd.n243 avdd.n242 1.83057
R1310 avdd.n244 avdd.n243 1.83057
R1311 avdd.n306 avdd.n0 1.72691
R1312 avdd.n241 avdd.n240 1.59141
R1313 avdd.n245 avdd.n240 1.59141
R1314 avdd.n228 avdd.n226 1.59141
R1315 avdd.n230 avdd.n228 1.59141
R1316 avdd.n252 avdd.n225 1.56301
R1317 avdd.n302 avdd.n301 1.33622
R1318 avdd.n206 avdd.n3 1.2505
R1319 avdd.n132 avdd.n94 1.2505
R1320 avdd.n166 avdd.n106 1.2505
R1321 avdd.n166 avdd.n165 1.2505
R1322 avdd.n167 avdd.n166 1.2505
R1323 avdd.n222 avdd.n5 1.2505
R1324 avdd.n222 avdd.n4 1.2505
R1325 avdd.n222 avdd.n221 1.2505
R1326 avdd.n238 avdd.n225 1.19516
R1327 avdd.n291 avdd.n252 1.01766
R1328 avdd.n301 avdd.n300 0.825743
R1329 avdd.n303 avdd.n225 0.691218
R1330 avdd.n2 avdd.n1 0.640571
R1331 avdd.n252 avdd.n251 0.5755
R1332 avdd.n268 avdd.n267 0.477136
R1333 avdd.n90 avdd.n2 0.466145
R1334 avdd.n149 avdd.n131 0.373307
R1335 avdd.n170 avdd.n126 0.373307
R1336 avdd.n181 avdd.n107 0.373307
R1337 avdd.n104 avdd.n95 0.373307
R1338 avdd.n205 avdd.n31 0.373307
R1339 avdd.n209 avdd.n7 0.373307
R1340 avdd.n218 avdd.n10 0.373307
R1341 avdd.n63 avdd.n62 0.373307
R1342 avdd.n304 avdd.n303 0.322423
R1343 avdd.n132 avdd.n3 0.283158
R1344 avdd.n224 avdd.n2 0.256667
R1345 avdd.n306 avdd.n305 0.222799
R1346 avdd.n305 avdd.n304 0.215455
R1347 avdd.n133 avdd.n132 0.173491
R1348 avdd.n278 avdd.n276 0.156463
R1349 avdd.n291 avdd.n290 0.141782
R1350 avdd.n223 avdd.n3 0.140453
R1351 avdd.n290 avdd.n289 0.138312
R1352 avdd.n303 avdd.n302 0.104705
R1353 avdd.n305 avdd.n1 0.0827949
R1354 avdd.n304 avdd.n224 0.0827949
R1355 avdd.n164 avdd.n126 0.0760556
R1356 avdd.n182 avdd.n181 0.0760556
R1357 avdd.n194 avdd.n95 0.0760556
R1358 avdd.n220 avdd.n7 0.0760556
R1359 avdd.n65 avdd.n10 0.0760556
R1360 avdd.n62 avdd.n60 0.0760556
R1361 avdd.n168 avdd.n131 0.0760556
R1362 avdd.n207 avdd.n205 0.0760556
R1363 avdd.n133 avdd.n1 0.06338
R1364 avdd.n224 avdd.n223 0.06338
R1365 avdd avdd.n306 0.0168616
R1366 avdd.n289 avdd 0.0161154
R1367 avdd.n290 avdd.n253 0.0043015
R1368 avdd.n302 avdd 0.0036996
R1369 avdd.n166 avdd.n133 0.000849819
R1370 avdd.n223 avdd.n222 0.000849819
R1371 dvdd.n18 dvdd.n13 1444.24
R1372 dvdd.n22 dvdd.n12 1444.24
R1373 dvdd.n22 dvdd.n13 1444.24
R1374 dvdd.n5 dvdd.n4 1444.24
R1375 dvdd.n26 dvdd.n25 1219.06
R1376 dvdd.n25 dvdd.n8 1219.06
R1377 dvdd.n37 dvdd.t2 954.721
R1378 dvdd.n0 dvdd.t4 941.715
R1379 dvdd.n6 dvdd.n5 774.586
R1380 dvdd.n34 dvdd.n3 766.821
R1381 dvdd.n31 dvdd.n3 656.23
R1382 dvdd.n31 dvdd.n6 648.687
R1383 dvdd.n26 dvdd.n6 547.413
R1384 dvdd.n8 dvdd.n3 547.413
R1385 dvdd.n24 dvdd.n23 491.368
R1386 dvdd.n32 dvdd.t3 474.889
R1387 dvdd.n24 dvdd.t3 471.904
R1388 dvdd.t5 dvdd.n32 471.904
R1389 dvdd.n23 dvdd.t0 375.529
R1390 dvdd.n33 dvdd.n4 365.901
R1391 dvdd.n39 dvdd.t6 324.887
R1392 dvdd.n9 dvdd.t1 324.589
R1393 dvdd.n18 dvdd.n17 317.007
R1394 dvdd.n20 dvdd.n19 181.986
R1395 dvdd.t5 dvdd.n5 159.195
R1396 dvdd.n20 dvdd.n12 143.627
R1397 dvdd.n16 dvdd.n13 140
R1398 dvdd.n13 dvdd.t0 140
R1399 dvdd.n27 dvdd.n26 140
R1400 dvdd.n26 dvdd.t3 140
R1401 dvdd.n35 dvdd.n34 140
R1402 dvdd.n28 dvdd.n5 140
R1403 dvdd.n14 dvdd.n8 140
R1404 dvdd.n8 dvdd.t3 140
R1405 dvdd.n19 dvdd.n16 132.814
R1406 dvdd.n28 dvdd.n2 120.847
R1407 dvdd.n34 dvdd.n33 103.171
R1408 dvdd.n29 dvdd.n28 99.7576
R1409 dvdd.n17 dvdd.n12 99.615
R1410 dvdd.n25 dvdd.n11 93.3338
R1411 dvdd.n25 dvdd.n24 93.3338
R1412 dvdd.n30 dvdd.n29 83.5434
R1413 dvdd.n30 dvdd.n1 76.2576
R1414 dvdd.n27 dvdd.n7 70.5005
R1415 dvdd.n29 dvdd.n27 70.5005
R1416 dvdd.n35 dvdd.n2 70.0696
R1417 dvdd.n19 dvdd.n18 70.0005
R1418 dvdd.n4 dvdd.n2 70.0005
R1419 dvdd.n31 dvdd.n30 70.0005
R1420 dvdd.n32 dvdd.n31 70.0005
R1421 dvdd.n22 dvdd.n21 70.0005
R1422 dvdd.n23 dvdd.n22 70.0005
R1423 dvdd.n21 dvdd.n20 58.6638
R1424 dvdd.n15 dvdd.n14 53.2047
R1425 dvdd.n33 dvdd.t5 38.7122
R1426 dvdd.n16 dvdd.n15 31.7338
R1427 dvdd.n17 dvdd.t0 30.7307
R1428 dvdd.n36 dvdd.n1 17.8809
R1429 dvdd.n14 dvdd.n1 16.5833
R1430 dvdd.n11 dvdd.n10 12.6415
R1431 dvdd.n37 dvdd.n36 5.7505
R1432 dvdd.n15 dvdd.n11 4.53383
R1433 dvdd.n10 dvdd.n9 3.83834
R1434 dvdd.n10 dvdd.n7 2.44153
R1435 dvdd.n21 dvdd.n7 0.610756
R1436 dvdd.n39 dvdd.n38 0.367833
R1437 dvdd.n40 dvdd.n39 0.178242
R1438 dvdd.n36 dvdd.n35 0.172217
R1439 dvdd.n40 dvdd.n0 0.169439
R1440 dvdd.n9 dvdd.n0 0.0715293
R1441 dvdd.n38 dvdd.n37 0.044
R1442 dvdd.n41 dvdd.n40 0.0263929
R1443 dvdd dvdd.n41 0.0263929
R1444 dvdd.n38 dvdd 0.005575
R1445 dvdd.n41 dvdd 0.001225
R1446 dvss.n42 dvss.n38 25476.2
R1447 dvss.n43 dvss.n19 9928.12
R1448 dvss.n62 dvss.n11 2461.06
R1449 dvss.n24 dvss.n11 2461.06
R1450 dvss.n62 dvss.n12 2461.06
R1451 dvss.n24 dvss.n12 2461.06
R1452 dvss.n40 dvss.n35 2125.76
R1453 dvss.n44 dvss.n35 2125.76
R1454 dvss.n44 dvss.n34 2125.76
R1455 dvss.n37 dvss.n9 2125.76
R1456 dvss.n65 dvss.n9 2125.76
R1457 dvss.n37 dvss.n10 2125.76
R1458 dvss.n65 dvss.n10 2125.76
R1459 dvss.n54 dvss.n22 2072.12
R1460 dvss.n22 dvss.n20 2072.12
R1461 dvss.n21 dvss.n20 2072.12
R1462 dvss.n54 dvss.n21 2072.12
R1463 dvss.n64 dvss.n63 1740.52
R1464 dvss.n56 dvss.n17 1629.53
R1465 dvss.n56 dvss.n18 1629.53
R1466 dvss.n49 dvss.n17 1629.53
R1467 dvss.n49 dvss.n18 1629.53
R1468 dvss.n25 dvss.n23 1449.84
R1469 dvss.n41 dvss.n40 862.641
R1470 dvss.n27 dvss.n26 850.245
R1471 dvss.t4 dvss.n43 818.846
R1472 dvss.n38 dvss.t2 667.819
R1473 dvss.n64 dvss.t2 667.819
R1474 dvss.n63 dvss.t6 569.837
R1475 dvss.n48 dvss.t5 468.853
R1476 dvss.n13 dvss.n11 422.277
R1477 dvss.n10 dvss.n8 420
R1478 dvss.t2 dvss.n10 420
R1479 dvss.n9 dvss.n7 420
R1480 dvss.t2 dvss.n9 420
R1481 dvss.n40 dvss.n39 420
R1482 dvss.n45 dvss.n44 420
R1483 dvss.n44 dvss.t4 420
R1484 dvss.n18 dvss.n15 420
R1485 dvss.t5 dvss.n18 420
R1486 dvss.n54 dvss.n53 420
R1487 dvss.t0 dvss.n54 420
R1488 dvss.n50 dvss.n49 420
R1489 dvss.n49 dvss.n48 420
R1490 dvss.n31 dvss.n17 420
R1491 dvss.t5 dvss.n17 420
R1492 dvss.n30 dvss.n20 420
R1493 dvss.t0 dvss.n20 420
R1494 dvss.n57 dvss.n56 420
R1495 dvss.n56 dvss.n55 420
R1496 dvss.n60 dvss.n12 420
R1497 dvss.n12 dvss.t6 420
R1498 dvss.n11 dvss.t6 420
R1499 dvss.n55 dvss.t0 367.87
R1500 dvss.n41 dvss.n34 365.515
R1501 dvss.n6 dvss.t1 357.413
R1502 dvss.n42 dvss.n41 351.276
R1503 dvss.n1 dvss.t3 341.531
R1504 dvss.n26 dvss.t6 317.377
R1505 dvss.n34 dvss.n33 280.243
R1506 dvss.n66 dvss.n65 280
R1507 dvss.n65 dvss.n64 280
R1508 dvss.n37 dvss.n36 280
R1509 dvss.n38 dvss.n37 280
R1510 dvss.n35 dvss.n32 280
R1511 dvss.n43 dvss.n35 280
R1512 dvss.n52 dvss.n22 280
R1513 dvss.n48 dvss.n22 280
R1514 dvss.n28 dvss.n21 280
R1515 dvss.n23 dvss.n21 280
R1516 dvss.n26 dvss.n25 252.459
R1517 dvss.t4 dvss.n42 233.216
R1518 dvss.n24 dvss.n14 210
R1519 dvss.n25 dvss.n24 210
R1520 dvss.n62 dvss.n61 210
R1521 dvss.n63 dvss.n62 210
R1522 dvss.n61 dvss.n60 183.5
R1523 dvss.n23 dvss.n19 155.083
R1524 dvss.n53 dvss.n52 154.732
R1525 dvss.n47 dvss.n46 134.024
R1526 dvss.n3 dvss.t7 124.424
R1527 dvss.n61 dvss.n13 115.001
R1528 dvss.n36 dvss.n8 114.392
R1529 dvss.n39 dvss.n33 108.769
R1530 dvss.t0 dvss.t5 100.984
R1531 dvss.n36 dvss.n7 99.4989
R1532 dvss.n45 dvss.n33 98.3464
R1533 dvss.n52 dvss.n51 75.7274
R1534 dvss.n58 dvss.n57 73.4648
R1535 dvss.n53 dvss.n29 70.5005
R1536 dvss.n60 dvss.n59 70.5005
R1537 dvss.n50 dvss.n47 63.9557
R1538 dvss.n39 dvss.n32 58.4049
R1539 dvss.n51 dvss.n50 56.7191
R1540 dvss.n66 dvss.n8 51.9346
R1541 dvss.n55 dvss.n19 46.8857
R1542 dvss.n30 dvss.n16 42.327
R1543 dvss.n57 dvss.n16 34.9112
R1544 dvss.n68 dvss.n67 22.8257
R1545 dvss.n46 dvss.n45 22.6667
R1546 dvss.n29 dvss.n6 21.0769
R1547 dvss.n68 dvss.n7 17.7561
R1548 dvss.n46 dvss.n32 16.1287
R1549 dvss.n27 dvss.n16 15.012
R1550 dvss.n59 dvss.n58 13.4258
R1551 dvss.n67 dvss.n1 11.5005
R1552 dvss.n51 dvss.n31 9.02218
R1553 dvss.n59 dvss.n14 8.77344
R1554 dvss.n58 dvss.n15 7.47521
R1555 dvss.n13 dvss.n2 7.438
R1556 dvss.n5 dvss.n0 6.743
R1557 dvss.n29 dvss.n28 6.31701
R1558 dvss.n70 dvss.n2 5.76655
R1559 dvss.n69 dvss.n68 4.17852
R1560 dvss.n67 dvss.n66 3.92358
R1561 dvss.n69 dvss.n6 3.63714
R1562 dvss.n3 dvss.n0 3.0455
R1563 dvss.n27 dvss.n2 2.50496
R1564 dvss.n31 dvss.n30 1.94336
R1565 dvss.n47 dvss.n15 1.45575
R1566 dvss.n4 dvss.n3 1.4505
R1567 dvss.n5 dvss 1.0155
R1568 dvss.n4 dvss 0.677167
R1569 dvss.n72 dvss.n0 0.508
R1570 dvss.n28 dvss.n27 0.351417
R1571 dvss.n69 dvss 0.138339
R1572 dvss.n70 dvss.n69 0.0892269
R1573 dvss.n16 dvss.n14 0.0784817
R1574 dvss.n71 dvss.n1 0.0622021
R1575 dvss.n70 dvss.n5 0.0547366
R1576 dvss.n71 dvss.n70 0.0153871
R1577 dvss.n72 dvss.n71 0.0144938
R1578 dvss.n5 dvss.n4 0.00216031
R1579 dvss dvss.n72 0.00198871
R1580 dvss.n4 dvss 0.00105343
R1581 dout.n1 dout.t0 362.913
R1582 dout.n0 dout.t2 343.055
R1583 dout.n0 dout.t1 324.56
R1584 dout.n1 dout.n0 8.50667
R1585 dout dout.n1 0.355381
C0 avss a_8004_3118# 0.273142f
C1 a_2174_9768# a_1842_9768# 0.321738f
C2 avdd a_700_3118# 0.322803f
C3 avss a_11304_7168# 0.185549f
C4 a_10162_518# avss 0.212389f
C5 a_8502_518# avss 0.212389f
C6 avdd a_8170_518# 0.013465f
C7 a_514_9768# avss 0.351175f
C8 avss a_700_3118# 1.41679f
C9 avdd a_9332_3118# 0.027973f
C10 avdd a_10992_3118# 0.010121f
C11 level_shifter_0.outb_h a_3082_4788# 0.212975f
C12 a_9146_9768# avdd 0.060792f
C13 avdd level_shifter_0.outb_h 2.10759f
C14 a_8170_518# avss 0.212389f
C15 dvdd level_shifter_0.out_h 0.036161f
C16 a_6344_3118# a_6012_3118# 0.321738f
C17 a_9810_9768# a_9478_9768# 0.321738f
C18 a_8834_518# a_9166_518# 0.321738f
C19 avss a_9332_3118# 0.246496f
C20 a_4684_3118# avss 0.36325f
C21 a_4020_3118# a_3688_3118# 0.321738f
C22 avdd a_680_7168# 0.04077f
C23 a_8170_518# a_7838_518# 0.321738f
C24 avdd a_7984_7168# 0.035787f
C25 avss a_10992_3118# 0.239858f
C26 level_shifter_0.outb_h avss 5.78953f
C27 avdd a_6086_5653# 1.21868f
C28 a_9146_9768# avss 0.181467f
C29 ena a_11636_7168# 0.16059f
C30 a_3668_7168# a_3336_7168# 0.321738f
C31 avss a_5680_3118# 1.43369f
C32 a_8980_7168# a_9312_7168# 0.321738f
C33 ena a_7560_4786# 0.179031f
C34 a_680_7168# avss 0.273825f
C35 a_7984_7168# avss 0.250638f
C36 level_shifter_0.out_h level_shifter_0.inb_l 0.32569f
C37 a_10660_3118# a_11636_7168# 0.016617f
C38 a_4020_3118# a_4352_3118# 0.321738f
C39 avdd a_1842_9768# 0.060792f
C40 avss a_6012_3118# 1.43369f
C41 a_2982_4700# a_5306_4788# 0.587047f
C42 a_6178_518# a_6510_518# 0.321738f
C43 avdd a_4750_4788# 1.65372f
C44 avdd a_1198_518# 0.013465f
C45 a_4036_4788# avss 1.20853f
C46 level_shifter_0.outb_h a_3638_4788# 0.219977f
C47 avss a_1842_9768# 0.181467f
C48 a_4664_7168# avdd 0.04474f
C49 dvdd a_11636_7168# 1.17978f
C50 avss a_4750_4788# 6.19241f
C51 avdd a_10142_9768# 0.060792f
C52 avss a_1198_518# 0.212389f
C53 a_5348_3118# a_5680_3118# 0.321738f
C54 a_2526_4188# avss 1.06716f
C55 avdd a_5660_7168# 1.20389f
C56 a_4664_7168# avss 0.250638f
C57 ena dvdd 2.35802f
C58 dout a_11636_7168# 0.117383f
C59 a_10142_9768# avss 0.181467f
C60 a_3834_9768# a_3502_9768# 0.321738f
C61 a_11324_3118# a_11636_7168# 0.337162f
C62 a_9146_9768# a_9478_9768# 0.321738f
C63 a_5660_7168# avss 0.250638f
C64 a_1414_4786# level_shifter_0.out_h 0.197567f
C65 ena dout 0.273692f
C66 a_11636_7168# level_shifter_0.inb_l 0.232978f
C67 a_10494_518# a_10162_518# 0.321738f
C68 a_4036_4788# a_3638_4788# 0.189325f
C69 a_6988_7168# a_7320_7168# 0.321738f
C70 level_shifter_0.outb_h a_6260_4788# 0.023308f
C71 a_2008_7168# avdd 0.048558f
C72 ena level_shifter_0.inb_l 1.19459f
C73 a_7008_3118# a_7340_3118# 0.321738f
C74 avdd a_1510_9768# 0.060792f
C75 a_4332_7168# avdd 0.051078f
C76 a_11158_518# a_11490_518# 0.321738f
C77 a_1032_3118# a_1364_3118# 0.321738f
C78 avdd a_3004_7168# 1.20389f
C79 a_2858_518# a_2526_518# 0.321738f
C80 avdd a_8714_4659# 0.567829f
C81 a_1414_4786# a_4194_4788# 0.011269f
C82 a_2008_7168# avss 0.250638f
C83 a_5862_4788# a_2982_4700# 0.671056f
C84 a_3854_518# avdd 0.013465f
C85 a_3356_3118# avss 1.22093f
C86 avss a_1510_9768# 0.181467f
C87 a_4332_7168# avss 0.250638f
C88 a_3006_5653# a_2982_4700# 0.120169f
C89 a_3004_7168# avss 0.250638f
C90 a_7008_3118# avss 0.795401f
C91 avss a_8714_4659# 0.041407f
C92 a_9000_3118# avdd 0.027973f
C93 avdd a_4854_5653# 0.98478f
C94 a_3854_518# avss 0.212389f
C95 a_514_7168# level_shifter_0.out_h 0.162381f
C96 dvdd dout 1.17946f
C97 level_shifter_0.out_h a_5306_4788# 0.350178f
C98 a_9000_3118# avss 0.24708f
C99 avdd a_8316_7168# 0.035899f
C100 a_2360_3118# a_2028_3118# 0.321738f
C101 dvdd level_shifter_0.inb_l 0.882379f
C102 a_3356_3118# a_3024_3118# 0.321738f
C103 a_8668_3118# avdd 0.027973f
C104 a_1012_7168# a_1344_7168# 0.321738f
C105 a_2368_4788# level_shifter_0.outb_h 0.088773f
C106 a_10660_3118# a_10328_3118# 0.321738f
C107 a_4592_4788# a_4194_4788# 0.188535f
C108 a_10328_3118# a_9996_3118# 0.321738f
C109 a_7154_9768# a_7486_9768# 0.321738f
C110 a_8004_3118# a_7672_3118# 0.321738f
C111 a_2982_4700# a_3082_4788# 0.972469f
C112 avss a_8316_7168# 0.27984f
C113 a_8502_518# a_8834_518# 0.321738f
C114 dout level_shifter_0.inb_l 0.189402f
C115 avdd a_2982_4700# 2.37155f
C116 a_8668_3118# avss 0.249073f
C117 a_9976_7168# a_9644_7168# 0.321738f
C118 a_1414_4786# a_5148_4788# 0.143491f
C119 avdd a_8336_3118# 0.027973f
C120 a_6086_5653# a_2368_4788# 0.145198f
C121 avdd a_3522_518# 0.013465f
C122 level_shifter_0.outb_h a_5704_4788# 0.023308f
C123 avdd a_9830_518# 0.013465f
C124 avss a_2982_4700# 5.56306f
C125 avdd a_7718_4786# 0.967771f
C126 a_1696_3118# a_1364_3118# 0.321738f
C127 a_8336_3118# avss 0.251575f
C128 avdd a_5328_7168# 0.933074f
C129 a_3522_518# avss 0.212389f
C130 avdd a_1862_518# 0.013465f
C131 avdd a_4996_7168# 0.054861f
C132 a_4194_4788# a_4238_5653# 0.017212f
C133 avdd a_846_9768# 0.060792f
C134 a_3622_5653# a_3082_4788# 0.128456f
C135 a_9830_518# avss 0.212389f
C136 avdd a_10474_9768# 0.060792f
C137 avdd a_3622_5653# 1.22095f
C138 a_7718_4786# avss 0.854394f
C139 a_2008_7168# a_2340_7168# 0.321738f
C140 a_2924_4788# level_shifter_0.outb_h 0.023308f
C141 a_6702_5653# a_2982_4700# 0.017212f
C142 a_8648_7168# a_8316_7168# 0.321738f
C143 avss a_5328_7168# 0.250638f
C144 avss a_1862_518# 0.212389f
C145 a_8502_518# a_8170_518# 0.321738f
C146 avdd a_4186_518# 0.013465f
C147 avss a_4996_7168# 0.250638f
C148 a_846_9768# avss 0.181467f
C149 a_3004_7168# a_3336_7168# 0.321738f
C150 a_2368_4788# a_4750_4788# 0.014269f
C151 avss a_10474_9768# 0.181467f
C152 level_shifter_0.out_h a_9482_5327# 0.120625f
C153 avdd a_5992_7168# 1.20389f
C154 a_2360_3118# a_2692_3118# 0.321738f
C155 a_2526_4188# a_2368_4788# 0.017212f
C156 level_shifter_0.out_h a_5862_4788# 0.3767f
C157 a_1178_9768# a_1510_9768# 0.321738f
C158 avss a_4186_518# 0.212389f
C159 a_3638_4788# a_2982_4700# 0.407234f
C160 a_5148_4788# a_5306_4788# 0.038465f
C161 avss a_5992_7168# 0.250638f
C162 a_10142_9768# a_9810_9768# 0.321738f
C163 avdd a_4000_7168# 0.780926f
C164 avdd a_2194_518# 0.013465f
C165 avdd a_2526_518# 0.013465f
C166 avss a_1364_3118# 0.299016f
C167 a_3622_5653# a_3638_4788# 0.047733f
C168 avdd a_9312_7168# 0.041727f
C169 a_1414_4786# a_3480_4788# 0.143491f
C170 a_2526_4188# a_2924_4788# 0.028806f
C171 a_6324_7168# a_5992_7168# 0.321738f
C172 avdd a_7652_7168# 0.041727f
C173 avdd a_6510_518# 0.013465f
C174 avss a_4000_7168# 0.250638f
C175 a_2174_9768# a_2506_9768# 0.321738f
C176 a_4518_518# a_4186_518# 0.321738f
C177 a_2194_518# avss 0.212389f
C178 level_shifter_0.out_h a_3082_4788# 0.409885f
C179 a_8814_9768# a_8482_9768# 0.321738f
C180 avss a_2526_518# 0.212389f
C181 avdd level_shifter_0.out_h 2.87832f
C182 a_6260_4788# a_2982_4700# 0.041881f
C183 avss a_9312_7168# 0.27984f
C184 a_3170_9768# a_3502_9768# 0.321738f
C185 a_7652_7168# avss 0.250638f
C186 a_7718_4786# a_11890_5939# 0.060633f
C187 avss a_6510_518# 0.212389f
C188 a_1012_7168# avdd 0.037216f
C189 a_6490_9768# avdd 0.060792f
C190 level_shifter_0.out_h avss 6.11633f
C191 avdd a_8814_9768# 0.060792f
C192 a_6012_3118# a_5680_3118# 0.321738f
C193 ena a_9482_5327# 0.117896f
C194 a_4036_4788# level_shifter_0.outb_h 0.023308f
C195 avdd a_4194_4788# 1.51515f
C196 a_2368_4788# a_4854_5653# 0.145198f
C197 a_1012_7168# avss 0.2747f
C198 a_6490_9768# avss 0.181467f
C199 a_5182_518# a_4850_518# 0.321738f
C200 level_shifter_0.outb_h a_4750_4788# 0.239282f
C201 a_8814_9768# avss 0.181467f
C202 a_1178_9768# a_846_9768# 0.321738f
C203 avdd a_6656_7168# 1.20389f
C204 a_9996_3118# a_9664_3118# 0.321738f
C205 a_2526_4188# level_shifter_0.outb_h 0.022591f
C206 a_4194_4788# avss 6.10201f
C207 a_5470_5653# a_5306_4788# 0.017212f
C208 avdd a_2672_7168# 1.20389f
C209 a_4020_3118# avss 0.42234f
C210 a_1696_3118# a_2028_3118# 0.321738f
C211 avss a_6656_7168# 0.250638f
C212 a_6490_9768# a_6158_9768# 0.321738f
C213 level_shifter_0.out_h a_3638_4788# 0.255355f
C214 avdd a_10972_7168# 1.26266f
C215 a_2368_4788# a_2982_4700# 0.011462f
C216 avdd a_11636_7168# 1.7381f
C217 avdd a_3502_9768# 0.060792f
C218 avdd a_2506_9768# 0.060792f
C219 a_2672_7168# avss 0.250638f
C220 avdd a_7560_4786# 0.023534f
C221 avdd a_9644_7168# 0.545447f
C222 a_1676_7168# a_1344_7168# 0.321738f
C223 avss a_10972_7168# 0.184602f
C224 ena avdd 2.33235f
C225 a_11636_7168# avss 0.998341f
C226 a_3502_9768# avss 0.181467f
C227 a_3522_518# a_3190_518# 0.321738f
C228 a_2506_9768# avss 0.181467f
C229 a_1414_4786# a_4592_4788# 0.143491f
C230 a_1414_4786# a_514_7168# 0.026766f
C231 a_3638_4788# a_4194_4788# 0.47078f
C232 avss a_7560_4786# 0.592294f
C233 a_6324_7168# a_6656_7168# 0.321738f
C234 a_9644_7168# avss 0.236063f
C235 a_2368_4788# a_3622_5653# 0.145198f
C236 a_10806_9768# avdd 0.060792f
C237 ena avss 1.46775f
C238 a_1414_4786# a_5306_4788# 0.011254f
C239 a_10660_3118# avdd 0.010121f
C240 avss a_5148_4788# 1.30325f
C241 avdd a_9996_3118# 0.015902f
C242 level_shifter_0.outb_h a_8714_4659# 0.30521f
C243 a_2924_4788# a_2982_4700# 0.171959f
C244 a_10806_9768# avss 0.181467f
C245 a_9000_3118# a_9332_3118# 0.321738f
C246 a_3688_3118# avss 0.378634f
C247 a_10660_3118# avss 0.239858f
C248 a_9996_3118# avss 0.239858f
C249 a_8336_3118# a_8004_3118# 0.321738f
C250 avss a_2028_3118# 1.43401f
C251 dvdd avdd 2.23594f
C252 a_10162_518# a_9830_518# 0.321738f
C253 avdd a_7486_9768# 0.060792f
C254 a_1842_9768# a_1510_9768# 0.321738f
C255 dout avdd 0.105337f
C256 avss a_4352_3118# 0.392067f
C257 dvdd avss 2.08884f
C258 a_3834_9768# avdd 0.060792f
C259 avdd a_9498_518# 0.013465f
C260 a_11324_3118# avdd 0.010121f
C261 a_7984_7168# a_8316_7168# 0.321738f
C262 a_7486_9768# avss 0.181467f
C263 a_6490_9768# a_6822_9768# 0.321738f
C264 a_2340_7168# a_2672_7168# 0.321738f
C265 avdd a_1530_518# 0.013465f
C266 a_514_9768# a_846_9768# 0.321738f
C267 a_3688_3118# a_3638_4788# 0.010379f
C268 level_shifter_0.outb_h a_2982_4700# 0.339321f
C269 avdd a_10826_518# 0.013465f
C270 a_6344_3118# a_6676_3118# 0.321738f
C271 a_7154_9768# avdd 0.060792f
C272 a_8980_7168# avdd 0.036775f
C273 avdd level_shifter_0.inb_l 0.591561f
C274 a_3668_7168# a_4000_7168# 0.321738f
C275 a_4332_7168# a_4664_7168# 0.321738f
C276 avdd a_4850_518# 0.013465f
C277 a_3834_9768# avss 0.181467f
C278 a_7652_7168# a_7320_7168# 0.321738f
C279 level_shifter_0.out_h a_2368_4788# 0.651754f
C280 a_9498_518# avss 0.212389f
C281 a_11324_3118# avss 0.239858f
C282 a_1414_4786# a_5862_4788# 0.011273f
C283 avss a_10826_518# 0.212389f
C284 a_3480_4788# a_3082_4788# 0.188913f
C285 a_1530_518# avss 0.212389f
C286 a_7718_4786# level_shifter_0.outb_h 0.257508f
C287 ena a_11890_5939# 0.287466f
C288 a_7154_9768# avss 0.181467f
C289 avdd a_5470_5653# 1.19052f
C290 level_shifter_0.inb_l avss 1.16675f
C291 a_4854_5653# a_4750_4788# 0.017212f
C292 a_8980_7168# avss 0.27984f
C293 avss a_4850_518# 0.212389f
C294 a_6842_518# a_6510_518# 0.321738f
C295 avdd a_6178_518# 0.013465f
C296 avdd a_11470_9768# 0.081826f
C297 avdd a_866_518# 0.013465f
C298 a_2360_3118# avss 1.43401f
C299 a_10640_7168# a_10972_7168# 0.321738f
C300 a_9976_7168# a_10308_7168# 0.321738f
C301 a_3480_4788# avss 1.2117f
C302 avss a_2692_3118# 1.43401f
C303 a_2368_4788# a_4194_4788# 0.016534f
C304 avdd a_10328_3118# 0.010421f
C305 a_6178_518# avss 0.212389f
C306 avss a_11470_9768# 0.352968f
C307 avss a_6676_3118# 1.43369f
C308 a_866_518# avss 0.212389f
C309 avdd a_1676_7168# 0.037821f
C310 a_7174_518# avdd 0.013465f
C311 a_10328_3118# avss 0.239858f
C312 a_9498_518# a_9166_518# 0.321738f
C313 a_2982_4700# a_4750_4788# 0.464544f
C314 a_8980_7168# a_8648_7168# 0.321738f
C315 a_8150_9768# a_8482_9768# 0.321738f
C316 a_1414_4786# a_3082_4788# 0.01694f
C317 a_1414_4786# avdd 0.013995f
C318 avss a_1676_7168# 0.266135f
C319 a_7174_518# avss 0.212389f
C320 a_2506_9768# a_2838_9768# 0.321738f
C321 a_4518_518# a_4850_518# 0.321738f
C322 dvdd a_11890_5939# 0.214298f
C323 a_3024_3118# a_2692_3118# 0.321738f
C324 a_7174_518# a_7506_518# 0.321738f
C325 a_5862_4788# a_5306_4788# 0.868266f
C326 a_4498_9768# a_4830_9768# 0.321738f
C327 a_3834_9768# a_4166_9768# 0.321738f
C328 avdd a_9976_7168# 1.26266f
C329 a_7818_9768# a_7486_9768# 0.321738f
C330 a_6988_7168# a_6656_7168# 0.321738f
C331 a_3480_4788# a_3638_4788# 0.038565f
C332 a_1414_4786# avss 15.251599f
C333 dout a_11890_5939# 0.799213f
C334 avdd a_8150_9768# 0.060792f
C335 a_4664_7168# a_4996_7168# 0.321738f
C336 a_9976_7168# avss 0.184602f
C337 a_8150_9768# avss 0.181467f
C338 a_5660_7168# a_5328_7168# 0.321738f
C339 a_10806_9768# a_11138_9768# 0.321738f
C340 a_10142_9768# a_10474_9768# 0.321738f
C341 level_shifter_0.out_h level_shifter_0.outb_h 4.31009f
C342 avdd a_2858_518# 0.013465f
C343 a_7652_7168# a_7984_7168# 0.321738f
C344 a_514_7168# avdd 0.76829f
C345 avdd a_1344_7168# 0.03676f
C346 a_5182_518# avdd 0.013465f
C347 a_2858_518# avss 0.212389f
C348 avdd a_5306_4788# 1.89931f
C349 a_9146_9768# a_8814_9768# 0.321738f
C350 a_4684_3118# a_4194_4788# 0.011588f
C351 a_8668_3118# a_9000_3118# 0.321738f
C352 a_1414_4786# a_3638_4788# 0.011114f
C353 a_1012_7168# a_680_7168# 0.321738f
C354 a_5660_7168# a_5992_7168# 0.321738f
C355 a_10972_7168# a_11304_7168# 0.321738f
C356 a_514_7168# avss 3.55411f
C357 a_4592_4788# avss 1.20861f
C358 a_6178_518# a_5846_518# 0.321738f
C359 level_shifter_0.outb_h a_4194_4788# 0.23346f
C360 a_11636_7168# a_11304_7168# 0.319467f
C361 a_3854_518# a_3522_518# 0.321738f
C362 a_10494_518# a_10826_518# 0.321738f
C363 a_1032_3118# avss 1.12081f
C364 a_4830_9768# avdd 0.060792f
C365 avss a_1344_7168# 0.2747f
C366 a_5182_518# avss 0.212389f
C367 avss a_5306_4788# 6.22238f
C368 a_7154_9768# a_6822_9768# 0.321738f
C369 avdd a_4238_5653# 1.00161f
C370 avdd a_5826_9768# 0.060792f
C371 a_4830_9768# avss 0.181467f
C372 a_4830_9768# a_5162_9768# 0.321738f
C373 a_6702_5653# a_5306_4788# 0.014515f
C374 level_shifter_0.out_h a_4750_4788# 0.324347f
C375 a_5826_9768# avss 0.181467f
C376 a_8668_3118# a_8336_3118# 0.321738f
C377 a_3854_518# a_4186_518# 0.321738f
C378 a_2526_4188# level_shifter_0.out_h 0.124112f
C379 a_5826_9768# a_5494_9768# 0.321738f
C380 a_11636_7168# a_10992_3118# 0.016617f
C381 a_1414_4786# a_6260_4788# 0.109899f
C382 a_4036_4788# a_4194_4788# 0.037969f
C383 a_7818_9768# a_8150_9768# 0.321738f
C384 level_shifter_0.outb_h a_7560_4786# 0.019812f
C385 a_2174_9768# avdd 0.060792f
C386 a_866_518# a_534_518# 0.321738f
C387 ena level_shifter_0.outb_h 0.572774f
C388 a_4194_4788# a_4750_4788# 0.504623f
C389 a_5470_5653# a_2368_4788# 0.145198f
C390 a_4498_9768# avdd 0.060792f
C391 a_11158_518# a_10826_518# 0.321738f
C392 avdd a_9664_3118# 0.02915f
C393 level_shifter_0.outb_h a_5148_4788# 0.023308f
C394 avdd a_3170_9768# 0.060792f
C395 avdd a_9482_5327# 0.683213f
C396 a_5826_9768# a_6158_9768# 0.321738f
C397 a_11138_9768# a_11470_9768# 0.321738f
C398 a_2174_9768# avss 0.181467f
C399 a_7718_4786# a_2982_4700# 0.247078f
C400 avdd a_5862_4788# 1.14612f
C401 a_5182_518# a_5514_518# 0.321738f
C402 a_4332_7168# a_4000_7168# 0.321738f
C403 a_10660_3118# a_10992_3118# 0.321738f
C404 a_4498_9768# avss 0.181467f
C405 a_9664_3118# avss 0.242783f
C406 a_3638_4788# a_4238_5653# 0.128681f
C407 a_3006_5653# a_3082_4788# 0.022867f
C408 a_3170_9768# avss 0.181467f
C409 avdd a_10308_7168# 1.26266f
C410 avdd a_3006_5653# 1.24299f
C411 a_1696_3118# avss 0.874205f
C412 a_5862_4788# avss 1.39834f
C413 avss a_5016_3118# 0.445627f
C414 a_4996_7168# a_5328_7168# 0.321738f
C415 avss a_10308_7168# 0.184602f
C416 level_shifter_0.out_h a_8714_4659# 0.405768f
C417 a_4684_3118# a_4352_3118# 0.321738f
C418 avdd a_8482_9768# 0.060792f
C419 a_6702_5653# a_5862_4788# 0.128965f
C420 dvdd level_shifter_0.outb_h 0.015481f
C421 a_6344_3118# avss 1.43369f
C422 a_6842_518# a_7174_518# 0.321738f
C423 a_5148_4788# a_4750_4788# 0.18926f
C424 avss a_8482_9768# 0.181467f
C425 avdd a_3082_4788# 1.75064f
C426 a_1414_4786# a_5704_4788# 0.143491f
C427 a_11324_3118# a_10992_3118# 0.321738f
C428 a_7340_3118# avss 0.403398f
C429 avss a_3082_4788# 5.91211f
C430 level_shifter_0.inb_l level_shifter_0.outb_h 0.26329f
C431 a_5348_3118# a_5016_3118# 0.321738f
C432 avdd avss 0.368908p
C433 a_4498_9768# a_4166_9768# 0.321738f
C434 avdd a_5494_9768# 0.060792f
C435 avdd a_7506_518# 0.013465f
C436 avdd a_5162_9768# 0.060792f
C437 a_4194_4788# a_4854_5653# 0.131849f
C438 a_1414_4786# a_2924_4788# 0.143491f
C439 avdd a_7838_518# 0.013465f
C440 a_3004_7168# a_2672_7168# 0.321738f
C441 a_514_7168# a_2368_4788# 0.099312f
C442 a_3480_4788# level_shifter_0.outb_h 0.023308f
C443 level_shifter_0.out_h a_2982_4700# 1.60036f
C444 avdd a_6702_5653# 1.22236f
C445 avss a_5494_9768# 0.181467f
C446 a_2194_518# a_1862_518# 0.321738f
C447 a_3190_518# a_2858_518# 0.321738f
C448 avss a_7506_518# 0.212389f
C449 avss a_5162_9768# 0.181467f
C450 a_5162_9768# a_5494_9768# 0.321738f
C451 avss a_7838_518# 0.212389f
C452 a_2368_4788# a_5306_4788# 0.015275f
C453 avdd a_6158_9768# 0.060792f
C454 a_7838_518# a_7506_518# 0.321738f
C455 a_6324_7168# avdd 1.20389f
C456 level_shifter_0.out_h a_7718_4786# 0.224983f
C457 avdd a_8648_7168# 0.035754f
C458 a_5862_4788# a_6260_4788# 0.203217f
C459 ena a_8714_4659# 0.049416f
C460 a_4194_4788# a_2982_4700# 0.365214f
C461 a_3638_4788# a_3082_4788# 0.753015f
C462 a_5704_4788# a_5306_4788# 0.194438f
C463 avdd a_9166_518# 0.013465f
C464 avdd a_3638_4788# 1.54584f
C465 avss a_6158_9768# 0.181467f
C466 avdd a_4518_518# 0.013465f
C467 a_2368_4788# a_4238_5653# 0.145198f
C468 a_3688_3118# a_3356_3118# 0.321738f
C469 a_6324_7168# avss 0.250638f
C470 a_3024_3118# avss 1.43401f
C471 a_1530_518# a_1198_518# 0.321738f
C472 a_8648_7168# avss 0.27984f
C473 avdd a_5514_518# 0.013465f
C474 avss a_9166_518# 0.212389f
C475 a_1414_4786# level_shifter_0.outb_h 0.179623f
C476 a_4518_518# avss 0.212389f
C477 a_3638_4788# avss 6.07746f
C478 avdd a_4166_9768# 0.060792f
C479 a_5348_3118# avss 1.33635f
C480 a_5470_5653# a_4750_4788# 0.134626f
C481 a_10640_7168# a_10308_7168# 0.321738f
C482 avdd a_9478_9768# 0.060792f
C483 avss a_5514_518# 0.212389f
C484 avdd a_7818_9768# 0.060792f
C485 avss a_4166_9768# 0.181467f
C486 a_3170_9768# a_2838_9768# 0.321738f
C487 a_866_518# a_1198_518# 0.321738f
C488 avdd a_5846_518# 0.013465f
C489 a_2194_518# a_2526_518# 0.321738f
C490 avdd a_3336_7168# 1.20389f
C491 avdd a_2340_7168# 0.823344f
C492 a_7560_4786# a_2982_4700# 0.228353f
C493 a_1032_3118# a_700_3118# 0.321738f
C494 avss a_9478_9768# 0.181467f
C495 a_7818_9768# avss 0.181467f
C496 ena a_2982_4700# 0.021677f
C497 a_1178_9768# avdd 0.060792f
C498 a_5862_4788# a_2368_4788# 0.013893f
C499 a_7718_4786# a_11636_7168# 0.104426f
C500 avss a_5846_518# 0.212389f
C501 a_3336_7168# avss 0.250638f
C502 a_2340_7168# avss 0.250638f
C503 a_1414_4786# a_4036_4788# 0.143491f
C504 a_7718_4786# a_7560_4786# 0.017316f
C505 avss a_6260_4788# 1.35888f
C506 a_4592_4788# level_shifter_0.outb_h 0.023308f
C507 a_514_7168# level_shifter_0.outb_h 0.111314f
C508 a_2368_4788# a_3006_5653# 0.145198f
C509 ena a_7718_4786# 0.649743f
C510 a_1178_9768# avss 0.181467f
C511 a_10640_7168# avdd 1.26266f
C512 a_1414_4786# a_4750_4788# 0.01122f
C513 a_10494_518# avdd 0.013465f
C514 a_5862_4788# a_5704_4788# 0.038138f
C515 level_shifter_0.outb_h a_5306_4788# 0.256952f
C516 a_514_7168# a_680_7168# 0.326105f
C517 level_shifter_0.inb_l a_8714_4659# 0.011544f
C518 a_1414_4786# a_2526_4188# 0.144624f
C519 avdd a_6822_9768# 0.060792f
C520 a_10640_7168# avss 0.184602f
C521 a_10494_518# avss 0.212389f
C522 avdd a_534_518# 0.034769f
C523 a_6086_5653# a_5306_4788# 0.139208f
C524 avdd a_2838_9768# 0.060792f
C525 a_10806_9768# a_10474_9768# 0.321738f
C526 avss a_6822_9768# 0.181467f
C527 dvdd a_2982_4700# 0.160393f
C528 level_shifter_0.out_h a_4194_4788# 0.29207f
C529 avdd a_11138_9768# 0.060792f
C530 a_2368_4788# a_3082_4788# 0.033098f
C531 a_7008_3118# a_6676_3118# 0.321738f
C532 avss a_534_518# 0.382983f
C533 avdd a_2368_4788# 13.213401f
C534 a_2008_7168# a_1676_7168# 0.321738f
C535 a_2838_9768# avss 0.181467f
C536 avdd a_7320_7168# 0.048021f
C537 avdd a_9810_9768# 0.060792f
C538 a_5846_518# a_5514_518# 0.321738f
C539 dvdd a_7718_4786# 1.46362f
C540 a_4592_4788# a_4750_4788# 0.03857f
C541 avss a_11138_9768# 0.181467f
C542 avdd a_3190_518# 0.013465f
C543 a_2368_4788# avss 0.50654f
C544 a_3668_7168# avdd 1.20389f
C545 a_11158_518# avdd 0.013465f
C546 a_7320_7168# avss 0.250638f
C547 a_6842_518# avdd 0.013465f
C548 a_4750_4788# a_5306_4788# 0.870813f
C549 a_9810_9768# avss 0.181467f
C550 dout a_7718_4786# 1.27607f
C551 avdd a_11490_518# 0.035085f
C552 a_9664_3118# a_9332_3118# 0.321738f
C553 a_6988_7168# avdd 0.663924f
C554 a_9830_518# a_9498_518# 0.321738f
C555 a_3190_518# avss 0.212389f
C556 a_9644_7168# a_9312_7168# 0.321738f
C557 a_3668_7168# avss 0.250638f
C558 avss a_5704_4788# 1.33621f
C559 a_11158_518# avss 0.212389f
C560 a_6702_5653# a_2368_4788# 0.145198f
C561 level_shifter_0.outb_h a_9482_5327# 0.221402f
C562 a_4684_3118# a_5016_3118# 0.321738f
C563 a_6842_518# avss 0.212389f
C564 a_8834_518# avdd 0.013465f
C565 a_2924_4788# a_3082_4788# 0.038253f
C566 a_11490_518# avss 0.382695f
C567 a_7340_3118# a_7672_3118# 0.321738f
C568 a_5862_4788# level_shifter_0.outb_h 0.2507f
C569 a_7718_4786# level_shifter_0.inb_l 1.00487f
C570 a_6988_7168# avss 0.250638f
C571 a_1530_518# a_1862_518# 0.321738f
C572 ena level_shifter_0.out_h 0.389292f
C573 avdd a_11304_7168# 1.08398f
C574 a_8834_518# avss 0.212389f
C575 a_6086_5653# a_5862_4788# 0.017212f
C576 a_2924_4788# avss 1.33599f
C577 a_2368_4788# a_3638_4788# 0.014219f
C578 avdd a_10162_518# 0.013465f
C579 a_8502_518# avdd 0.013465f
C580 avss a_7672_3118# 0.310838f
C581 a_514_9768# avdd 0.082099f
C582 dout dvss 1.76453f
C583 ena dvss 2.512052f
C584 dvdd dvss 9.599436f
C585 avss dvss 6.051995f
C586 avdd dvss 0.393525p
C587 a_11490_518# dvss 0.392297f
C588 a_11324_3118# dvss 0.340341f
C589 a_11158_518# dvss 0.358381f
C590 a_10992_3118# dvss 0.340341f
C591 a_10826_518# dvss 0.358381f
C592 a_10660_3118# dvss 0.340341f
C593 a_10494_518# dvss 0.358381f
C594 a_10328_3118# dvss 0.352273f
C595 a_10162_518# dvss 0.358381f
C596 a_9996_3118# dvss 0.353394f
C597 a_9830_518# dvss 0.358381f
C598 a_9664_3118# dvss 0.340341f
C599 a_9498_518# dvss 0.358381f
C600 a_9332_3118# dvss 0.340341f
C601 a_9166_518# dvss 0.358381f
C602 a_9000_3118# dvss 0.340341f
C603 a_8834_518# dvss 0.358381f
C604 a_8668_3118# dvss 0.340341f
C605 a_8502_518# dvss 0.358381f
C606 a_8336_3118# dvss 0.340341f
C607 a_8170_518# dvss 0.358381f
C608 a_8004_3118# dvss 0.340341f
C609 a_7838_518# dvss 0.358381f
C610 a_7672_3118# dvss 0.340341f
C611 a_7506_518# dvss 0.358381f
C612 a_7340_3118# dvss 0.340341f
C613 a_7174_518# dvss 0.358381f
C614 a_7008_3118# dvss 0.340341f
C615 a_6842_518# dvss 0.358381f
C616 a_6676_3118# dvss 0.340341f
C617 a_6510_518# dvss 0.358381f
C618 a_6344_3118# dvss 0.340341f
C619 a_6178_518# dvss 0.358381f
C620 a_6012_3118# dvss 0.340341f
C621 a_5846_518# dvss 0.358381f
C622 a_5680_3118# dvss 0.340341f
C623 a_5514_518# dvss 0.358381f
C624 a_5348_3118# dvss 0.340341f
C625 a_5182_518# dvss 0.358381f
C626 a_5016_3118# dvss 0.340341f
C627 a_4850_518# dvss 0.358381f
C628 a_4684_3118# dvss 0.340341f
C629 a_4518_518# dvss 0.358381f
C630 a_4352_3118# dvss 0.340341f
C631 a_4186_518# dvss 0.358381f
C632 a_4020_3118# dvss 0.340341f
C633 a_3854_518# dvss 0.358381f
C634 a_3688_3118# dvss 0.340341f
C635 a_3522_518# dvss 0.358381f
C636 a_3356_3118# dvss 0.340341f
C637 a_3190_518# dvss 0.358381f
C638 a_3024_3118# dvss 0.340341f
C639 a_2858_518# dvss 0.358381f
C640 a_2692_3118# dvss 0.340341f
C641 a_2526_518# dvss 0.358381f
C642 a_2360_3118# dvss 0.340341f
C643 a_2194_518# dvss 0.358381f
C644 a_2028_3118# dvss 0.340341f
C645 a_1862_518# dvss 0.358381f
C646 a_1696_3118# dvss 0.340341f
C647 a_1530_518# dvss 0.358381f
C648 a_1364_3118# dvss 0.340341f
C649 a_1198_518# dvss 0.358381f
C650 a_1032_3118# dvss 0.34253f
C651 a_866_518# dvss 0.358381f
C652 a_700_3118# dvss 0.346799f
C653 a_534_518# dvss 0.391326f
C654 a_11890_5939# dvss 0.814248f
C655 a_7560_4786# dvss 0.0144f
C656 a_6260_4788# dvss 0.012204f
C657 a_5704_4788# dvss 0.012204f
C658 a_5148_4788# dvss 0.012204f
C659 a_4592_4788# dvss 0.012204f
C660 a_4036_4788# dvss 0.012204f
C661 a_3480_4788# dvss 0.012204f
C662 a_2924_4788# dvss 0.014421f
C663 a_2526_4188# dvss 0.012204f
C664 a_1414_4786# dvss 0.764141f
C665 a_9482_5327# dvss 0.011184f
C666 a_8714_4659# dvss 0.010821f
C667 level_shifter_0.outb_h dvss 0.480526f
C668 level_shifter_0.inb_l dvss 1.27748f
C669 a_7718_4786# dvss 1.12939f
C670 a_5862_4788# dvss 0.175811f
C671 a_5306_4788# dvss 0.400428f
C672 a_4750_4788# dvss 0.314033f
C673 a_4194_4788# dvss 0.326912f
C674 a_3638_4788# dvss 0.31549f
C675 a_3082_4788# dvss 0.459116f
C676 a_2982_4700# dvss 0.489027f
C677 level_shifter_0.out_h dvss 0.629318f
C678 a_6702_5653# dvss 0.011305f
C679 a_6086_5653# dvss 0.011305f
C680 a_5470_5653# dvss 0.011305f
C681 a_4854_5653# dvss 0.011305f
C682 a_4238_5653# dvss 0.011305f
C683 a_3622_5653# dvss 0.011305f
C684 a_3006_5653# dvss 0.011305f
C685 a_2368_4788# dvss 0.677014f
C686 a_11636_7168# dvss 3.97595f
C687 a_11470_9768# dvss 0.391386f
C688 a_11304_7168# dvss 0.338939f
C689 a_11138_9768# dvss 0.358545f
C690 a_10972_7168# dvss 0.338762f
C691 a_10806_9768# dvss 0.358545f
C692 a_10640_7168# dvss 0.338762f
C693 a_10474_9768# dvss 0.358545f
C694 a_10308_7168# dvss 0.338762f
C695 a_10142_9768# dvss 0.358545f
C696 a_9976_7168# dvss 0.338762f
C697 a_9810_9768# dvss 0.358545f
C698 a_9644_7168# dvss 0.340651f
C699 a_9478_9768# dvss 0.358545f
C700 a_9312_7168# dvss 0.338762f
C701 a_9146_9768# dvss 0.358545f
C702 a_8980_7168# dvss 0.338762f
C703 a_8814_9768# dvss 0.358545f
C704 a_8648_7168# dvss 0.338762f
C705 a_8482_9768# dvss 0.358545f
C706 a_8316_7168# dvss 0.338762f
C707 a_8150_9768# dvss 0.358545f
C708 a_7984_7168# dvss 0.338762f
C709 a_7818_9768# dvss 0.358545f
C710 a_7652_7168# dvss 0.338762f
C711 a_7486_9768# dvss 0.358545f
C712 a_7320_7168# dvss 0.338762f
C713 a_7154_9768# dvss 0.358545f
C714 a_6988_7168# dvss 0.338762f
C715 a_6822_9768# dvss 0.358545f
C716 a_6656_7168# dvss 0.338762f
C717 a_6490_9768# dvss 0.358545f
C718 a_6324_7168# dvss 0.338762f
C719 a_6158_9768# dvss 0.358545f
C720 a_5992_7168# dvss 0.338762f
C721 a_5826_9768# dvss 0.358545f
C722 a_5660_7168# dvss 0.338762f
C723 a_5494_9768# dvss 0.358545f
C724 a_5328_7168# dvss 0.338762f
C725 a_5162_9768# dvss 0.358545f
C726 a_4996_7168# dvss 0.338762f
C727 a_4830_9768# dvss 0.358545f
C728 a_4664_7168# dvss 0.338762f
C729 a_4498_9768# dvss 0.358545f
C730 a_4332_7168# dvss 0.338762f
C731 a_4166_9768# dvss 0.358545f
C732 a_4000_7168# dvss 0.338762f
C733 a_3834_9768# dvss 0.358545f
C734 a_3668_7168# dvss 0.338762f
C735 a_3502_9768# dvss 0.358545f
C736 a_3336_7168# dvss 0.338762f
C737 a_3170_9768# dvss 0.358545f
C738 a_3004_7168# dvss 0.338762f
C739 a_2838_9768# dvss 0.358545f
C740 a_2672_7168# dvss 0.338762f
C741 a_2506_9768# dvss 0.358545f
C742 a_2340_7168# dvss 0.338762f
C743 a_2174_9768# dvss 0.358545f
C744 a_2008_7168# dvss 0.338762f
C745 a_1842_9768# dvss 0.358545f
C746 a_1676_7168# dvss 0.338762f
C747 a_1510_9768# dvss 0.358545f
C748 a_1344_7168# dvss 0.338762f
C749 a_1178_9768# dvss 0.358545f
C750 a_1012_7168# dvss 0.338762f
C751 a_846_9768# dvss 0.358545f
C752 a_680_7168# dvss 0.338762f
C753 a_514_7168# dvss 0.18866f
C754 a_514_9768# dvss 0.392573f
C755 dvdd.t4 dvss 0.010971f
C756 dvdd.n0 dvss 0.111155f
C757 dvdd.t2 dvss 0.020105f
C758 dvdd.n1 dvss 0.060181f
C759 dvdd.n2 dvss 0.075625f
C760 dvdd.n3 dvss 0.021959f
C761 dvdd.n4 dvss 0.153814f
C762 dvdd.n5 dvss 0.030763f
C763 dvdd.t3 dvss 0.169281f
C764 dvdd.n6 dvss 0.021946f
C765 dvdd.n7 dvss 0.013726f
C766 dvdd.n8 dvss 0.018955f
C767 dvdd.t1 dvss 0.025914f
C768 dvdd.n9 dvss 0.166731f
C769 dvdd.n10 dvss 0.039918f
C770 dvdd.n11 dvss 0.045384f
C771 dvdd.t0 dvss 0.239889f
C772 dvdd.n12 dvss 0.031614f
C773 dvdd.n13 dvss 0.031457f
C774 dvdd.n14 dvss 0.089105f
C775 dvdd.n15 dvss 0.055728f
C776 dvdd.n16 dvss 0.044651f
C777 dvdd.n18 dvss 0.18037f
C778 dvdd.n19 dvss 0.030189f
C779 dvdd.n20 dvss 0.076658f
C780 dvdd.n21 dvss 0.084672f
C781 dvdd.n22 dvss 0.031046f
C782 dvdd.n23 dvss 0.201093f
C783 dvdd.n24 dvss 0.161958f
C784 dvdd.n25 dvss 0.026601f
C785 dvdd.n26 dvss 0.018955f
C786 dvdd.n27 dvss 0.011328f
C787 dvdd.n28 dvss 0.026499f
C788 dvdd.n29 dvss 0.021946f
C789 dvdd.n30 dvss 0.013603f
C790 dvdd.n31 dvss 0.014307f
C791 dvdd.n32 dvss 0.169281f
C792 dvdd.t5 dvss 0.2913f
C793 dvdd.n34 dvss 0.028532f
C794 dvdd.n35 dvss 0.073843f
C795 dvdd.n36 dvss 0.036799f
C796 dvdd.n37 dvss 1.82245f
C797 dvdd.n38 dvss 0.016505f
C798 dvdd.t6 dvss 0.025959f
C799 dvdd.n39 dvss 0.062162f
C800 dvdd.n40 dvss 0.129417f
C801 dvdd.n41 dvss 0.132557f
C802 avdd.n0 dvss 14.0698f
C803 avdd.n1 dvss 6.83284f
C804 avdd.n2 dvss 4.06185f
C805 avdd.n3 dvss 0.708527f
C806 avdd.t1 dvss 0.022647f
C807 avdd.n4 dvss 0.480934f
C808 avdd.t3 dvss 0.022647f
C809 avdd.n5 dvss 0.480934f
C810 avdd.t11 dvss 0.022647f
C811 avdd.n6 dvss 0.042406f
C812 avdd.n7 dvss 0.14127f
C813 avdd.n8 dvss 0.036668f
C814 avdd.n9 dvss 0.037496f
C815 avdd.n10 dvss 0.14127f
C816 avdd.n11 dvss 0.129096f
C817 avdd.n12 dvss 0.129019f
C818 avdd.n13 dvss 0.129019f
C819 avdd.n14 dvss 1.33038f
C820 avdd.n15 dvss 0.129096f
C821 avdd.n16 dvss 1.33038f
C822 avdd.n17 dvss 0.129019f
C823 avdd.n18 dvss 0.129019f
C824 avdd.n19 dvss 0.174203f
C825 avdd.n20 dvss 0.174203f
C826 avdd.n21 dvss 0.129019f
C827 avdd.n22 dvss 0.129019f
C828 avdd.n23 dvss 1.33038f
C829 avdd.n24 dvss 0.129096f
C830 avdd.n25 dvss 0.129096f
C831 avdd.n26 dvss 1.33038f
C832 avdd.n27 dvss 0.036668f
C833 avdd.n28 dvss 0.129019f
C834 avdd.n29 dvss 0.037496f
C835 avdd.n30 dvss 0.042406f
C836 avdd.n31 dvss 0.121004f
C837 avdd.n32 dvss 0.129019f
C838 avdd.n33 dvss 0.043226f
C839 avdd.n34 dvss 0.043226f
C840 avdd.n35 dvss 0.037496f
C841 avdd.n36 dvss 0.273019f
C842 avdd.n37 dvss 0.129019f
C843 avdd.n38 dvss 0.129019f
C844 avdd.n39 dvss 2.16888f
C845 avdd.n40 dvss 0.129096f
C846 avdd.n41 dvss 1.33038f
C847 avdd.n42 dvss 0.129096f
C848 avdd.n43 dvss 0.129019f
C849 avdd.n44 dvss 0.129019f
C850 avdd.n45 dvss 0.549759f
C851 avdd.n46 dvss 0.037496f
C852 avdd.n47 dvss 1.22796f
C853 avdd.n48 dvss 1.18147f
C854 avdd.n49 dvss 0.129019f
C855 avdd.n50 dvss 0.348105f
C856 avdd.n51 dvss 0.273019f
C857 avdd.n52 dvss 0.302545f
C858 avdd.n53 dvss 0.129096f
C859 avdd.n55 dvss 2.16635f
C860 avdd.t23 dvss 1.68252f
C861 avdd.n56 dvss 0.129096f
C862 avdd.n57 dvss 0.143848f
C863 avdd.n58 dvss 0.372123f
C864 avdd.n59 dvss 0.042406f
C865 avdd.n60 dvss 0.373175f
C866 avdd.n61 dvss 0.043226f
C867 avdd.n62 dvss 0.14127f
C868 avdd.n63 dvss 0.121004f
C869 avdd.n64 dvss 0.042406f
C870 avdd.n65 dvss 0.233395f
C871 avdd.n66 dvss 0.25084f
C872 avdd.n67 dvss 0.036668f
C873 avdd.n68 dvss 0.174203f
C874 avdd.n69 dvss 0.164894f
C875 avdd.n70 dvss 0.129096f
C876 avdd.t2 dvss 1.4063f
C877 avdd.n71 dvss 0.129096f
C878 avdd.n72 dvss 0.164894f
C879 avdd.n73 dvss 0.1747f
C880 avdd.n74 dvss 0.1747f
C881 avdd.n75 dvss 0.164894f
C882 avdd.n76 dvss 0.1747f
C883 avdd.n77 dvss 0.1747f
C884 avdd.n78 dvss 0.164894f
C885 avdd.n79 dvss 0.1747f
C886 avdd.n80 dvss 0.1747f
C887 avdd.n81 dvss 0.129096f
C888 avdd.n82 dvss 0.129096f
C889 avdd.t12 dvss 1.4063f
C890 avdd.n83 dvss 0.129096f
C891 avdd.n84 dvss 0.036668f
C892 avdd.n85 dvss 0.129019f
C893 avdd.n86 dvss 0.129019f
C894 avdd.t4 dvss 1.4063f
C895 avdd.n87 dvss 0.129096f
C896 avdd.n88 dvss 0.129096f
C897 avdd.n89 dvss 0.14401f
C898 avdd.n90 dvss 2.02762f
C899 avdd.n91 dvss 0.112639f
C900 avdd.n92 dvss 0.174203f
C901 avdd.n93 dvss 0.174203f
C902 avdd.t5 dvss 0.022647f
C903 avdd.n94 dvss 0.480934f
C904 avdd.n95 dvss 0.14127f
C905 avdd.n96 dvss 0.164894f
C906 avdd.n97 dvss 0.043226f
C907 avdd.n98 dvss 0.1747f
C908 avdd.n99 dvss 0.129096f
C909 avdd.n100 dvss 0.037496f
C910 avdd.n101 dvss 1.33038f
C911 avdd.n102 dvss 0.164894f
C912 avdd.n103 dvss 0.174203f
C913 avdd.n104 dvss 0.121004f
C914 avdd.n105 dvss 0.042406f
C915 avdd.t9 dvss 0.022647f
C916 avdd.n106 dvss 0.480934f
C917 avdd.n107 dvss 0.121004f
C918 avdd.n108 dvss 0.1747f
C919 avdd.n109 dvss 0.129096f
C920 avdd.n110 dvss 0.129019f
C921 avdd.n111 dvss 0.164894f
C922 avdd.n112 dvss 1.33038f
C923 avdd.n113 dvss 0.129096f
C924 avdd.n114 dvss 0.129019f
C925 avdd.n115 dvss 0.129019f
C926 avdd.n116 dvss 0.174203f
C927 avdd.n117 dvss 0.036668f
C928 avdd.n118 dvss 0.042406f
C929 avdd.n119 dvss 0.174203f
C930 avdd.n120 dvss 0.129019f
C931 avdd.n121 dvss 0.129019f
C932 avdd.n122 dvss 1.33038f
C933 avdd.n123 dvss 0.129096f
C934 avdd.n124 dvss 0.129096f
C935 avdd.n125 dvss 1.33038f
C936 avdd.n126 dvss 0.14127f
C937 avdd.n127 dvss 0.036668f
C938 avdd.n128 dvss 0.129019f
C939 avdd.n129 dvss 0.037496f
C940 avdd.n130 dvss 0.042406f
C941 avdd.n131 dvss 0.14127f
C942 avdd.t15 dvss 0.022647f
C943 avdd.n132 dvss 0.763917f
C944 avdd.n133 dvss 2.71291f
C945 avdd.t7 dvss 0.022647f
C946 avdd.n134 dvss 0.129019f
C947 avdd.n135 dvss 0.043226f
C948 avdd.n136 dvss 0.043226f
C949 avdd.n137 dvss 0.28285f
C950 avdd.n138 dvss 0.129019f
C951 avdd.n139 dvss 0.129019f
C952 avdd.n140 dvss 1.33038f
C953 avdd.n141 dvss 0.129096f
C954 avdd.n142 dvss 1.33038f
C955 avdd.n143 dvss 0.129096f
C956 avdd.n144 dvss 0.129019f
C957 avdd.n145 dvss 0.129019f
C958 avdd.n146 dvss 0.174203f
C959 avdd.n147 dvss 0.128615f
C960 avdd.n148 dvss 0.089843f
C961 avdd.n149 dvss 0.145427f
C962 avdd.n150 dvss 0.30851f
C963 avdd.n151 dvss 0.088367f
C964 avdd.n152 dvss 0.280039f
C965 avdd.n153 dvss 0.271001f
C966 avdd.n154 dvss 0.129096f
C967 avdd.t14 dvss 1.4063f
C968 avdd.n155 dvss 0.129096f
C969 avdd.n156 dvss 0.272918f
C970 avdd.n157 dvss 0.1747f
C971 avdd.n158 dvss 0.1747f
C972 avdd.n159 dvss 0.164894f
C973 avdd.n160 dvss 0.1747f
C974 avdd.n161 dvss 0.1747f
C975 avdd.n162 dvss 0.037496f
C976 avdd.n163 dvss 0.25084f
C977 avdd.n164 dvss 0.233395f
C978 avdd.n165 dvss 0.480934f
C979 avdd.n166 dvss 1.25936f
C980 avdd.t22 dvss 0.022658f
C981 avdd.n167 dvss 0.645829f
C982 avdd.n168 dvss 0.233395f
C983 avdd.n169 dvss 0.25084f
C984 avdd.n170 dvss 0.121004f
C985 avdd.n171 dvss 0.129096f
C986 avdd.t6 dvss 1.4063f
C987 avdd.n172 dvss 0.129096f
C988 avdd.n173 dvss 0.164894f
C989 avdd.n174 dvss 0.174203f
C990 avdd.n175 dvss 0.174203f
C991 avdd.n176 dvss 0.164894f
C992 avdd.n177 dvss 0.129096f
C993 avdd.t8 dvss 1.4063f
C994 avdd.n178 dvss 0.129096f
C995 avdd.n179 dvss 0.129019f
C996 avdd.n180 dvss 0.043226f
C997 avdd.n181 dvss 0.14127f
C998 avdd.n182 dvss 0.233395f
C999 avdd.n183 dvss 0.25084f
C1000 avdd.n184 dvss 0.036668f
C1001 avdd.n185 dvss 0.129019f
C1002 avdd.n186 dvss 1.33038f
C1003 avdd.n187 dvss 0.129019f
C1004 avdd.n188 dvss 0.129096f
C1005 avdd.n189 dvss 0.164894f
C1006 avdd.n190 dvss 0.1747f
C1007 avdd.n191 dvss 0.1747f
C1008 avdd.n192 dvss 0.037496f
C1009 avdd.n193 dvss 0.25084f
C1010 avdd.n194 dvss 0.233395f
C1011 avdd.n195 dvss 0.042406f
C1012 avdd.n196 dvss 0.129019f
C1013 avdd.n197 dvss 1.33038f
C1014 avdd.n198 dvss 1.33038f
C1015 avdd.n199 dvss 0.129019f
C1016 avdd.n200 dvss 0.129096f
C1017 avdd.n201 dvss 0.129019f
C1018 avdd.n202 dvss 1.33038f
C1019 avdd.n203 dvss 0.129019f
C1020 avdd.n204 dvss 0.043226f
C1021 avdd.n205 dvss 0.14127f
C1022 avdd.t13 dvss 0.022647f
C1023 avdd.n206 dvss 0.480934f
C1024 avdd.n207 dvss 0.233395f
C1025 avdd.n208 dvss 0.25084f
C1026 avdd.n209 dvss 0.121004f
C1027 avdd.n210 dvss 0.129096f
C1028 avdd.t10 dvss 1.4063f
C1029 avdd.n211 dvss 0.129096f
C1030 avdd.n212 dvss 0.164894f
C1031 avdd.n213 dvss 0.174203f
C1032 avdd.n214 dvss 0.174203f
C1033 avdd.n215 dvss 0.164894f
C1034 avdd.n216 dvss 0.129096f
C1035 avdd.t0 dvss 1.4063f
C1036 avdd.n217 dvss 0.129096f
C1037 avdd.n218 dvss 0.121004f
C1038 avdd.n219 dvss 0.25084f
C1039 avdd.n220 dvss 0.233395f
C1040 avdd.n221 dvss 0.480934f
C1041 avdd.n222 dvss 1.25936f
C1042 avdd.n223 dvss 3.00063f
C1043 avdd.n224 dvss 5.98315f
C1044 avdd.n225 dvss 2.59915f
C1045 avdd.n226 dvss 6.58312f
C1046 avdd.n227 dvss 1.19324f
C1047 avdd.n228 dvss 3.4539f
C1048 avdd.n229 dvss 0.990578f
C1049 avdd.n230 dvss 14.805901f
C1050 avdd.n231 dvss 3.259f
C1051 avdd.n232 dvss 1.7832f
C1052 avdd.n233 dvss 0.814121f
C1053 avdd.n234 dvss 0.129096f
C1054 avdd.n235 dvss 0.129096f
C1055 avdd.n236 dvss 0.339033f
C1056 avdd.n237 dvss 0.144037f
C1057 avdd.n238 dvss 1.03799f
C1058 avdd.n239 dvss 2.72402f
C1059 avdd.n240 dvss 3.45408f
C1060 avdd.n241 dvss 4.90067f
C1061 avdd.n242 dvss 3.50538f
C1062 avdd.n243 dvss 4.05907f
C1063 avdd.n244 dvss 17.519499f
C1064 avdd.n245 dvss 14.8067f
C1065 avdd.n246 dvss 8.44591f
C1066 avdd.n247 dvss 1.9707f
C1067 avdd.n248 dvss 0.9904f
C1068 avdd.n249 dvss 1.64593f
C1069 avdd.n250 dvss 0.936816f
C1070 avdd.n251 dvss 0.807219f
C1071 avdd.n252 dvss 1.46402f
C1072 avdd.t17 dvss 0.022626f
C1073 avdd.n253 dvss 0.282641f
C1074 avdd.t20 dvss 0.022626f
C1075 avdd.n254 dvss 0.135889f
C1076 avdd.n255 dvss 0.258486f
C1077 avdd.n256 dvss 0.129019f
C1078 avdd.n257 dvss 0.129019f
C1079 avdd.n258 dvss 1.5174f
C1080 avdd.n259 dvss 0.129096f
C1081 avdd.n260 dvss 0.129096f
C1082 avdd.n261 dvss 1.54033f
C1083 avdd.n262 dvss 0.621898f
C1084 avdd.n263 dvss 0.196993f
C1085 avdd.n264 dvss 0.129096f
C1086 avdd.n265 dvss 0.235881f
C1087 avdd.n266 dvss 0.129019f
C1088 avdd.n267 dvss 0.135456f
C1089 avdd.n268 dvss 0.102113f
C1090 avdd.n269 dvss 0.129096f
C1091 avdd.t16 dvss 0.814121f
C1092 avdd.t21 dvss 0.814121f
C1093 avdd.n270 dvss 0.156509f
C1094 avdd.n271 dvss 0.26612f
C1095 avdd.n272 dvss 0.129019f
C1096 avdd.n273 dvss 0.814121f
C1097 avdd.n274 dvss 0.726211f
C1098 avdd.n275 dvss 0.129019f
C1099 avdd.n276 dvss 0.121004f
C1100 avdd.n277 dvss 0.129019f
C1101 avdd.n278 dvss 0.148071f
C1102 avdd.n279 dvss 0.307395f
C1103 avdd.n280 dvss 0.19446f
C1104 avdd.n281 dvss 0.129019f
C1105 avdd.n282 dvss 0.228632f
C1106 avdd.n283 dvss 0.337509f
C1107 avdd.n284 dvss 0.235056f
C1108 avdd.n285 dvss 0.129096f
C1109 avdd.t18 dvss 1.62224f
C1110 avdd.n286 dvss 0.129096f
C1111 avdd.n287 dvss 0.147507f
C1112 avdd.n288 dvss 0.173126f
C1113 avdd.n289 dvss -0.077995f
C1114 avdd.n290 dvss -2.3234f
C1115 avdd.n291 dvss 1.82343f
C1116 avdd.n292 dvss 0.175531f
C1117 avdd.n293 dvss 0.139614f
C1118 avdd.n294 dvss 0.129019f
C1119 avdd.n295 dvss 1.08549f
C1120 avdd.n296 dvss 4.34889f
C1121 avdd.n297 dvss 4.04848f
C1122 avdd.n298 dvss 8.4489f
C1123 avdd.n299 dvss 1.97142f
C1124 avdd.n300 dvss 0.693642f
C1125 avdd.n301 dvss 2.63538f
C1126 avdd.n302 dvss 7.82406f
C1127 avdd.n303 dvss 34.713898f
C1128 avdd.n304 dvss 39.6382f
C1129 avdd.n305 dvss 32.987698f
C1130 avdd.n306 dvss 22.104f
C1131 ena.t3 dvss 0.048434f
C1132 ena.t2 dvss 0.049086f
C1133 ena.t5 dvss 0.03596f
C1134 ena.t6 dvss 0.036608f
C1135 ena.n0 dvss 0.397742f
C1136 ena.n1 dvss 0.46328f
C1137 ena.t1 dvss 0.177359f
C1138 ena.t0 dvss 0.19358f
C1139 ena.n2 dvss 1.86542f
C1140 ena.t4 dvss 0.056172f
C1141 ena.n3 dvss 0.34841f
C1142 ena.n4 dvss 0.332895f
C1143 ena.n5 dvss 0.387439f
C1144 avss.n0 dvss 6.88022f
C1145 avss.n1 dvss 1.53256f
C1146 avss.n2 dvss 2.16361f
C1147 avss.n3 dvss 0.651011f
C1148 avss.n4 dvss 0.651011f
C1149 avss.t115 dvss 0.690506f
C1150 avss.n5 dvss 0.067816f
C1151 avss.n6 dvss 0.067816f
C1152 avss.n7 dvss 0.163153f
C1153 avss.n8 dvss 0.079751f
C1154 avss.t30 dvss 0.012228f
C1155 avss.n9 dvss 0.26078f
C1156 avss.n10 dvss 0.153856f
C1157 avss.n11 dvss 2.27039f
C1158 avss.n12 dvss 11.4207f
C1159 avss.t9 dvss 0.012133f
C1160 avss.n13 dvss 0.073914f
C1161 avss.n14 dvss 0.019321f
C1162 avss.n15 dvss 0.019321f
C1163 avss.n16 dvss 0.019366f
C1164 avss.n17 dvss 0.019321f
C1165 avss.n18 dvss 0.067816f
C1166 avss.t5 dvss 0.012134f
C1167 avss.n19 dvss 0.19429f
C1168 avss.n20 dvss 0.045077f
C1169 avss.n21 dvss 0.067963f
C1170 avss.n22 dvss 0.067963f
C1171 avss.t47 dvss 1.40074f
C1172 avss.n23 dvss 0.067816f
C1173 avss.t59 dvss 1.24291f
C1174 avss.n24 dvss 0.081266f
C1175 avss.n25 dvss 0.019366f
C1176 avss.n26 dvss 0.081896f
C1177 avss.t122 dvss 1.24949f
C1178 avss.n27 dvss 1.01274f
C1179 avss.t81 dvss 1.39312f
C1180 avss.n28 dvss 0.651011f
C1181 avss.n29 dvss 0.651011f
C1182 avss.n30 dvss 2.16199f
C1183 avss.n31 dvss 2.0716f
C1184 avss.n32 dvss 0.402545f
C1185 avss.t75 dvss 0.012113f
C1186 avss.n33 dvss 0.224131f
C1187 avss.n34 dvss 0.34155f
C1188 avss.n35 dvss 0.444186f
C1189 avss.n36 dvss 2.08339f
C1190 avss.t111 dvss 1.54459f
C1191 avss.t159 dvss 1.48764f
C1192 avss.t154 dvss 1.48764f
C1193 avss.t148 dvss 1.48764f
C1194 avss.t68 dvss 1.48764f
C1195 avss.t57 dvss 1.48764f
C1196 avss.t49 dvss 1.48764f
C1197 avss.t92 dvss 1.48764f
C1198 avss.t25 dvss 1.48764f
C1199 avss.t42 dvss 1.48764f
C1200 avss.t105 dvss 1.48764f
C1201 avss.t91 dvss 1.48974f
C1202 avss.t116 dvss 1.60193f
C1203 avss.t108 dvss 1.59997f
C1204 avss.t157 dvss 1.59997f
C1205 avss.t141 dvss 1.59997f
C1206 avss.t112 dvss 1.46021f
C1207 avss.t55 dvss 1.6004f
C1208 avss.t28 dvss 1.6004f
C1209 avss.t89 dvss 1.6004f
C1210 avss.t155 dvss 1.6004f
C1211 avss.t52 dvss 1.6004f
C1212 avss.t71 dvss 1.6004f
C1213 avss.t94 dvss 1.6004f
C1214 avss.t40 dvss 1.6004f
C1215 avss.t37 dvss 1.6004f
C1216 avss.t102 dvss 1.6004f
C1217 avss.t160 dvss 1.6004f
C1218 avss.t143 dvss 1.6004f
C1219 avss.t32 dvss 1.6004f
C1220 avss.t106 dvss 1.6004f
C1221 avss.t88 dvss 1.6004f
C1222 avss.t64 dvss 1.6004f
C1223 avss.t22 dvss 1.6004f
C1224 avss.t117 dvss 1.6004f
C1225 avss.t87 dvss 1.6004f
C1226 avss.t46 dvss 1.6004f
C1227 avss.t45 dvss 1.6004f
C1228 avss.t60 dvss 1.6004f
C1229 avss.t50 dvss 1.6004f
C1230 avss.t82 dvss 1.6004f
C1231 avss.t33 dvss 1.6004f
C1232 avss.t163 dvss 1.6004f
C1233 avss.t126 dvss 1.6004f
C1234 avss.t79 dvss 1.2003f
C1235 avss.n37 dvss 0.800202f
C1236 avss.t101 dvss 1.2003f
C1237 avss.t107 dvss 1.6004f
C1238 avss.t72 dvss 1.6004f
C1239 avss.t140 dvss 1.6004f
C1240 avss.t96 dvss 1.6004f
C1241 avss.t34 dvss 1.60042f
C1242 avss.t146 dvss 1.59999f
C1243 avss.t97 dvss 1.59997f
C1244 avss.t150 dvss 1.59997f
C1245 avss.t26 dvss 1.59997f
C1246 avss.t76 dvss 1.59997f
C1247 avss.t145 dvss 1.59997f
C1248 avss.t134 dvss 1.59997f
C1249 avss.t139 dvss 1.59997f
C1250 avss.t86 dvss 1.59997f
C1251 avss.t118 dvss 1.59997f
C1252 avss.t78 dvss 0.93974f
C1253 avss.n38 dvss 1.07907f
C1254 avss.n39 dvss 0.067816f
C1255 avss.n40 dvss 0.067816f
C1256 avss.n41 dvss 0.065747f
C1257 avss.n42 dvss 0.100546f
C1258 avss.n43 dvss 0.171545f
C1259 avss.n44 dvss 0.581921f
C1260 avss.n45 dvss 0.067963f
C1261 avss.t100 dvss 0.012142f
C1262 avss.n46 dvss 1.00752f
C1263 avss.n47 dvss 0.11676f
C1264 avss.t74 dvss 0.349845f
C1265 avss.t35 dvss 1.83067f
C1266 avss.n48 dvss 0.067982f
C1267 avss.t80 dvss 1.14427f
C1268 avss.n49 dvss 0.067816f
C1269 avss.n50 dvss 0.067816f
C1270 avss.n51 dvss 0.148277f
C1271 avss.n52 dvss 0.019277f
C1272 avss.n53 dvss 0.5922f
C1273 avss.n54 dvss 0.067963f
C1274 avss.t132 dvss 1.34813f
C1275 avss.n55 dvss 0.067816f
C1276 avss.n56 dvss 0.067963f
C1277 avss.t149 dvss 1.3284f
C1278 avss.n57 dvss 0.067816f
C1279 avss.n58 dvss 0.067816f
C1280 avss.n59 dvss 0.019321f
C1281 avss.n60 dvss 0.865492f
C1282 avss.n61 dvss 0.084953f
C1283 avss.n62 dvss 0.067816f
C1284 avss.n63 dvss 0.063944f
C1285 avss.t131 dvss 0.012913f
C1286 avss.n64 dvss 0.381025f
C1287 avss.n65 dvss 0.742642f
C1288 avss.t15 dvss 0.012133f
C1289 avss.n66 dvss 0.073914f
C1290 avss.n67 dvss 0.019321f
C1291 avss.n68 dvss 0.019321f
C1292 avss.n69 dvss 0.019321f
C1293 avss.n70 dvss 0.019321f
C1294 avss.n71 dvss 0.067816f
C1295 avss.n72 dvss 0.045634f
C1296 avss.n73 dvss 0.067963f
C1297 avss.n74 dvss 0.067963f
C1298 avss.t153 dvss 1.40074f
C1299 avss.n75 dvss 0.067816f
C1300 avss.t142 dvss 1.34813f
C1301 avss.n76 dvss 0.080882f
C1302 avss.n77 dvss 0.019321f
C1303 avss.n78 dvss 0.019321f
C1304 avss.n79 dvss 0.080882f
C1305 avss.n80 dvss 0.067963f
C1306 avss.n81 dvss 0.067963f
C1307 avss.t147 dvss 1.21661f
C1308 avss.n82 dvss 0.067816f
C1309 avss.n83 dvss 0.067816f
C1310 avss.t109 dvss 1.40074f
C1311 avss.n84 dvss 0.092224f
C1312 avss.n85 dvss 0.019321f
C1313 avss.n86 dvss 0.063944f
C1314 avss.t17 dvss 0.012133f
C1315 avss.n87 dvss 0.193424f
C1316 avss.n88 dvss 0.31838f
C1317 avss.n89 dvss 0.343743f
C1318 avss.t3 dvss 0.012133f
C1319 avss.n90 dvss 0.073914f
C1320 avss.n91 dvss 0.019321f
C1321 avss.n92 dvss 0.019321f
C1322 avss.n93 dvss 0.019321f
C1323 avss.n94 dvss 0.019321f
C1324 avss.n95 dvss 0.067816f
C1325 avss.n96 dvss 0.045634f
C1326 avss.n97 dvss 0.067963f
C1327 avss.n98 dvss 0.067963f
C1328 avss.t123 dvss 1.40074f
C1329 avss.n99 dvss 0.067816f
C1330 avss.t66 dvss 1.29552f
C1331 avss.n100 dvss 0.080882f
C1332 avss.n101 dvss 0.019321f
C1333 avss.n102 dvss 0.019321f
C1334 avss.n103 dvss 0.080882f
C1335 avss.n104 dvss 0.067963f
C1336 avss.n105 dvss 0.067963f
C1337 avss.t83 dvss 1.26922f
C1338 avss.n106 dvss 0.067816f
C1339 avss.n107 dvss 0.067816f
C1340 avss.t73 dvss 1.40074f
C1341 avss.n108 dvss 0.092224f
C1342 avss.n109 dvss 0.019321f
C1343 avss.n110 dvss 0.019321f
C1344 avss.n111 dvss 0.019321f
C1345 avss.n112 dvss 0.019321f
C1346 avss.n113 dvss 0.063944f
C1347 avss.t61 dvss 1.19688f
C1348 avss.n114 dvss 0.067963f
C1349 avss.t166 dvss 1.22318f
C1350 avss.n115 dvss 0.986438f
C1351 avss.n116 dvss 0.960133f
C1352 avss.n117 dvss 0.067963f
C1353 avss.n118 dvss 0.019321f
C1354 avss.n119 dvss 0.080882f
C1355 avss.n120 dvss 0.067963f
C1356 avss.n121 dvss 0.067963f
C1357 avss.t120 dvss 1.40074f
C1358 avss.n122 dvss 0.067816f
C1359 avss.t77 dvss 1.40074f
C1360 avss.n123 dvss 0.067816f
C1361 avss.n124 dvss 0.019321f
C1362 avss.n125 dvss 0.063944f
C1363 avss.t54 dvss 1.14427f
C1364 avss.n126 dvss 0.067963f
C1365 avss.t43 dvss 1.27579f
C1366 avss.n127 dvss 1.03905f
C1367 avss.n128 dvss 0.907523f
C1368 avss.n129 dvss 0.067963f
C1369 avss.n130 dvss 0.019321f
C1370 avss.n131 dvss 0.080882f
C1371 avss.n132 dvss 0.067963f
C1372 avss.n133 dvss 0.067963f
C1373 avss.t84 dvss 1.40074f
C1374 avss.n134 dvss 0.067816f
C1375 avss.t85 dvss 1.40074f
C1376 avss.n135 dvss 0.067816f
C1377 avss.n136 dvss 0.067963f
C1378 avss.n137 dvss 0.067963f
C1379 avss.n138 dvss 1.09166f
C1380 avss.t119 dvss 0.854913f
C1381 avss.n139 dvss 1.09166f
C1382 avss.n140 dvss 0.067963f
C1383 avss.n141 dvss 0.019321f
C1384 avss.n142 dvss 0.092224f
C1385 avss.n143 dvss 0.019321f
C1386 avss.t41 dvss 1.40074f
C1387 avss.t63 dvss 1.164f
C1388 avss.t18 dvss 1.09166f
C1389 avss.n144 dvss 0.067816f
C1390 avss.n145 dvss 0.136233f
C1391 avss.n146 dvss 0.145147f
C1392 avss.n147 dvss 0.23533f
C1393 avss.n148 dvss 0.23542f
C1394 avss.n149 dvss 0.088483f
C1395 avss.n150 dvss 0.080882f
C1396 avss.n151 dvss 0.019321f
C1397 avss.n152 dvss 0.067963f
C1398 avss.n153 dvss 1.09166f
C1399 avss.t48 dvss 0.690506f
C1400 avss.n154 dvss 0.710235f
C1401 avss.n155 dvss 0.545829f
C1402 avss.n156 dvss 0.067963f
C1403 avss.n157 dvss 0.019321f
C1404 avss.n158 dvss 0.080882f
C1405 avss.n159 dvss 0.080882f
C1406 avss.n160 dvss 0.080882f
C1407 avss.n161 dvss 0.088483f
C1408 avss.n162 dvss 0.067816f
C1409 avss.t14 dvss 1.09166f
C1410 avss.n163 dvss 0.067816f
C1411 avss.n164 dvss 0.088483f
C1412 avss.n165 dvss 0.080882f
C1413 avss.n166 dvss 0.080882f
C1414 avss.n167 dvss 0.088483f
C1415 avss.n168 dvss 0.080882f
C1416 avss.n169 dvss 0.080882f
C1417 avss.n170 dvss 0.08163f
C1418 avss.n171 dvss 2.76239f
C1419 avss.n172 dvss 1.06781f
C1420 avss.n173 dvss 0.043494f
C1421 avss.n174 dvss 0.019321f
C1422 avss.n175 dvss 0.067963f
C1423 avss.n176 dvss 1.09166f
C1424 avss.t144 dvss 0.854913f
C1425 avss.n177 dvss 1.09166f
C1426 avss.n178 dvss 0.067963f
C1427 avss.n179 dvss 0.067963f
C1428 avss.n180 dvss 1.09166f
C1429 avss.t24 dvss 0.854913f
C1430 avss.n181 dvss 1.09166f
C1431 avss.n182 dvss 0.067963f
C1432 avss.n183 dvss 0.019321f
C1433 avss.n184 dvss 0.092224f
C1434 avss.n185 dvss 0.019321f
C1435 avss.n186 dvss 0.080882f
C1436 avss.n187 dvss 0.080882f
C1437 avss.n188 dvss 0.088483f
C1438 avss.n189 dvss 0.067816f
C1439 avss.t2 dvss 1.09166f
C1440 avss.n190 dvss 0.067816f
C1441 avss.n191 dvss 0.088483f
C1442 avss.n192 dvss 0.080882f
C1443 avss.n193 dvss 0.080882f
C1444 avss.n194 dvss 0.088483f
C1445 avss.n195 dvss 0.080882f
C1446 avss.n196 dvss 0.080882f
C1447 avss.n197 dvss 0.088483f
C1448 avss.n198 dvss 0.080882f
C1449 avss.n199 dvss 0.080882f
C1450 avss.n200 dvss 0.067816f
C1451 avss.n201 dvss 0.063644f
C1452 avss.n202 dvss 0.067963f
C1453 avss.n203 dvss 0.07018f
C1454 avss.n204 dvss 0.330789f
C1455 avss.n205 dvss 0.080882f
C1456 avss.n206 dvss 0.080882f
C1457 avss.n207 dvss 0.088483f
C1458 avss.n208 dvss 0.067816f
C1459 avss.n209 dvss 0.067963f
C1460 avss.n210 dvss 1.09166f
C1461 avss.t128 dvss 0.854913f
C1462 avss.t0 dvss 1.40074f
C1463 avss.n211 dvss 0.080882f
C1464 avss.n212 dvss 0.080865f
C1465 avss.n213 dvss 0.088483f
C1466 avss.n214 dvss 0.067816f
C1467 avss.n215 dvss 0.067963f
C1468 avss.n216 dvss 0.067963f
C1469 avss.n217 dvss 0.067963f
C1470 avss.n218 dvss 1.09166f
C1471 avss.t51 dvss 0.854913f
C1472 avss.n219 dvss 1.09166f
C1473 avss.t103 dvss 1.40074f
C1474 avss.t8 dvss 1.09166f
C1475 avss.n220 dvss 0.067816f
C1476 avss.n221 dvss 0.067963f
C1477 avss.n222 dvss 1.09166f
C1478 avss.n223 dvss 0.067963f
C1479 avss.n224 dvss 0.019321f
C1480 avss.n225 dvss 0.092224f
C1481 avss.n226 dvss 0.063944f
C1482 avss.t13 dvss 0.012133f
C1483 avss.n227 dvss 0.193424f
C1484 avss.n228 dvss 1.28134f
C1485 avss.n229 dvss 0.687754f
C1486 avss.n230 dvss 1.581f
C1487 avss.t7 dvss 0.012133f
C1488 avss.n231 dvss 0.193424f
C1489 avss.n232 dvss 0.045634f
C1490 avss.n233 dvss 0.073914f
C1491 avss.n234 dvss 0.067816f
C1492 avss.t6 dvss 1.09166f
C1493 avss.n235 dvss 0.067816f
C1494 avss.n236 dvss 0.088483f
C1495 avss.n237 dvss 0.080882f
C1496 avss.n238 dvss 0.080882f
C1497 avss.n239 dvss 0.088483f
C1498 avss.n240 dvss 0.067816f
C1499 avss.t12 dvss 1.09166f
C1500 avss.n241 dvss 0.067816f
C1501 avss.n242 dvss 0.073914f
C1502 avss.n243 dvss 0.092224f
C1503 avss.n244 dvss 0.063944f
C1504 avss.n245 dvss 0.045634f
C1505 avss.n246 dvss 0.193424f
C1506 avss.n247 dvss 0.41346f
C1507 avss.n248 dvss 0.438709f
C1508 avss.t11 dvss 0.012133f
C1509 avss.n249 dvss 0.193424f
C1510 avss.n250 dvss 0.045634f
C1511 avss.n251 dvss 0.073914f
C1512 avss.n252 dvss 0.067816f
C1513 avss.t10 dvss 1.09166f
C1514 avss.n253 dvss 0.067816f
C1515 avss.n254 dvss 0.088483f
C1516 avss.n255 dvss 0.080882f
C1517 avss.n256 dvss 0.080882f
C1518 avss.n257 dvss 0.088483f
C1519 avss.n258 dvss 0.067816f
C1520 avss.t16 dvss 1.09166f
C1521 avss.n259 dvss 0.067816f
C1522 avss.n260 dvss 0.073914f
C1523 avss.n261 dvss 0.092224f
C1524 avss.n262 dvss 0.063944f
C1525 avss.n263 dvss 0.045634f
C1526 avss.n264 dvss 0.193424f
C1527 avss.n265 dvss 1.7112f
C1528 avss.n266 dvss 1.33669f
C1529 avss.n267 dvss 0.656076f
C1530 avss.n268 dvss 1.54043f
C1531 avss.t67 dvss 1.89613f
C1532 avss.t151 dvss 1.65505f
C1533 avss.t70 dvss 1.65505f
C1534 avss.t124 dvss 1.65505f
C1535 avss.t156 dvss 1.65505f
C1536 avss.t27 dvss 1.65505f
C1537 avss.t130 dvss 1.65505f
C1538 avss.t104 dvss 1.64635f
C1539 avss.t165 dvss 1.48034f
C1540 avss.t69 dvss 1.4859f
C1541 avss.t133 dvss 1.4859f
C1542 avss.t113 dvss 1.4859f
C1543 avss.t129 dvss 1.4859f
C1544 avss.t152 dvss 1.4859f
C1545 avss.t121 dvss 1.4859f
C1546 avss.t93 dvss 1.4859f
C1547 avss.t158 dvss 1.4859f
C1548 avss.t95 dvss 1.4859f
C1549 avss.t137 dvss 1.4859f
C1550 avss.t58 dvss 1.52695f
C1551 avss.n269 dvss 1.91853f
C1552 avss.n270 dvss 1.19741f
C1553 avss.n271 dvss 1.51883f
C1554 avss.n272 dvss 15.2899f
C1555 avss.n273 dvss 2.32651f
C1556 avss.t164 dvss 3.30636f
C1557 avss.n274 dvss 1.66678f
C1558 avss.t110 dvss 2.4194f
C1559 avss.n275 dvss 2.1338f
C1560 avss.t31 dvss 1.78251f
C1561 avss.n276 dvss 2.13361f
C1562 avss.t36 dvss 1.78251f
C1563 avss.t44 dvss 2.10691f
C1564 avss.n277 dvss 2.1716f
C1565 avss.n278 dvss 1.79166f
C1566 avss.n279 dvss 0.385744f
C1567 avss.n280 dvss 9.1536f
C1568 avss.n281 dvss 17.268301f
C1569 avss.n282 dvss 2.74237f
C1570 avss.t19 dvss 0.012133f
C1571 avss.n283 dvss 0.193424f
C1572 avss.n284 dvss 0.045634f
C1573 avss.n285 dvss 0.070272f
C1574 avss.n286 dvss 0.099537f
C1575 avss.n287 dvss 0.316653f
C1576 avss.n288 dvss 0.067963f
C1577 avss.n289 dvss 1.09166f
C1578 avss.t161 dvss 1.94657f
C1579 avss.t1 dvss 2.18332f
C1580 avss.t127 dvss 2.18332f
C1581 avss.t56 dvss 2.18332f
C1582 avss.t20 dvss 1.61776f
C1583 avss.n290 dvss 0.067963f
C1584 avss.n291 dvss 1.09166f
C1585 avss.t90 dvss 1.40074f
C1586 avss.t98 dvss 1.09166f
C1587 avss.n292 dvss 0.067816f
C1588 avss.n293 dvss 0.090923f
C1589 avss.n294 dvss 0.109565f
C1590 avss.n295 dvss 0.15829f
C1591 avss.n296 dvss 0.149315f
C1592 avss.n297 dvss 0.067963f
C1593 avss.n298 dvss 1.09166f
C1594 avss.t138 dvss 2.13071f
C1595 avss.t39 dvss 1.39417f
C1596 avss.n299 dvss 1.8233f
C1597 avss.n300 dvss 1.66656f
C1598 avss.n301 dvss 0.067963f
C1599 avss.n302 dvss 0.172753f
C1600 avss.n303 dvss 0.117195f
C1601 avss.n304 dvss 0.044673f
C1602 avss.n305 dvss 0.083242f
C1603 avss.n306 dvss 0.149475f
C1604 avss.n307 dvss 0.046407f
C1605 avss.n308 dvss 0.067816f
C1606 avss.t99 dvss 0.647549f
C1607 avss.n310 dvss 0.067816f
C1608 avss.n311 dvss 0.101164f
C1609 avss.n312 dvss 0.158692f
C1610 avss.n313 dvss 0.075341f
C1611 avss.n314 dvss 0.067963f
C1612 avss.n315 dvss 0.27909f
C1613 avss.n316 dvss 0.103576f
C1614 avss.n317 dvss 3.14054f
C1615 avss.n318 dvss 0.113274f
C1616 avss.n319 dvss 1.08706f
C1617 avss.n320 dvss 2.77268f
C1618 avss.n321 dvss 6.01835f
C1619 avss.n322 dvss 1.98945f
C1620 avss.t21 dvss 1.65195f
C1621 avss.t136 dvss 1.6004f
C1622 avss.t65 dvss 1.6004f
C1623 avss.t53 dvss 1.6004f
C1624 avss.t135 dvss 1.00748f
C1625 avss.n323 dvss 4.10924f
C1626 avss.n324 dvss 4.17053f
C1627 avss.t29 dvss 0.940404f
C1628 avss.t162 dvss 1.32183f
C1629 avss.t114 dvss 1.17057f
C1630 avss.n325 dvss 0.933828f
C1631 avss.n326 dvss 0.067963f
C1632 avss.n327 dvss 0.019366f
C1633 avss.n328 dvss 0.081251f
C1634 avss.n329 dvss 0.081251f
C1635 avss.n330 dvss 0.089042f
C1636 avss.n331 dvss 0.067816f
C1637 avss.t4 dvss 1.09166f
C1638 avss.n332 dvss 0.067816f
C1639 avss.n333 dvss 0.073013f
C1640 avss.n334 dvss 0.091547f
C1641 avss.n335 dvss 0.063975f
C1642 avss.n336 dvss 0.045634f
C1643 avss.n337 dvss 0.193424f
C1644 avss.n338 dvss 1.71327f
C1645 avss.n339 dvss 1.21878f
C1646 avss.n340 dvss 1.97282f
C1647 avss.n341 dvss 6.9573f
C1648 avss.n342 dvss 0.241842f
C1649 avss.n343 dvss 0.146961f
C1650 avss.n344 dvss 0.128004f
C1651 avss.n345 dvss 0.179153f
C1652 avss.n346 dvss 0.067963f
C1653 avss.n347 dvss 1.09166f
C1654 avss.t23 dvss 1.64406f
C1655 avss.t125 dvss 2.18332f
C1656 avss.t62 dvss 2.18332f
C1657 avss.t38 dvss 2.34641f
C1658 avss.n348 dvss 2.64662f
C1659 avss.n349 dvss 1.21372f
C1660 avss.n350 dvss 0.911706f
C1661 avss.n351 dvss 1.89424f
.ends

