magic
tech sky130A
magscale 1 2
timestamp 1699547976
<< dnwell >>
rect 116 6766 12126 10608
rect 116 3954 9974 6766
rect 116 116 12126 3954
<< nwell >>
rect 0 10402 12242 10724
rect 0 322 322 10402
rect 11920 6972 12242 10402
rect 7118 6034 7988 6713
rect 9768 6650 12242 6972
rect 7118 5356 7372 6034
rect 9768 4070 10090 6650
rect 11613 5041 11667 5393
rect 9768 3748 12242 4070
rect 11920 322 12242 3748
rect 0 0 12242 322
<< mvnsubdiff >>
rect 73 10631 12169 10651
rect 73 10597 153 10631
rect 12089 10597 12169 10631
rect 73 10577 12169 10597
rect 73 10571 147 10577
rect 73 153 93 10571
rect 127 153 147 10571
rect 12095 10571 12169 10577
rect 12095 6817 12115 10571
rect 12149 6817 12169 10571
rect 12095 6797 12169 6817
rect 9943 6777 12169 6797
rect 9943 6743 10048 6777
rect 12079 6743 12169 6777
rect 9943 6723 12169 6743
rect 9943 6695 10017 6723
rect 9943 4029 9963 6695
rect 9997 4029 10017 6695
rect 9943 3997 10017 4029
rect 9943 3977 12169 3997
rect 9943 3943 10048 3977
rect 12078 3943 12169 3977
rect 9943 3923 12169 3943
rect 73 147 147 153
rect 12095 3909 12169 3923
rect 12095 153 12115 3909
rect 12149 153 12169 3909
rect 12095 147 12169 153
rect 73 127 12169 147
rect 73 93 153 127
rect 12089 93 12169 127
rect 73 73 12169 93
<< mvnsubdiffcont >>
rect 153 10597 12089 10631
rect 93 153 127 10571
rect 12115 6817 12149 10571
rect 10048 6743 12079 6777
rect 9963 4029 9997 6695
rect 10048 3943 12078 3977
rect 12115 153 12149 3909
rect 153 93 12089 127
<< locali >>
rect 86 10631 12151 10636
rect 86 10597 153 10631
rect 12089 10597 12151 10631
rect 86 10571 12151 10597
rect 86 153 93 10571
rect 127 10493 12115 10571
rect 127 7683 210 10493
rect 193 4005 210 7683
rect 295 10295 11944 10409
rect 295 7090 409 10295
rect 11830 7090 11944 10295
rect 295 7071 11944 7090
rect 295 6986 8302 7071
rect 9743 6986 11944 7071
rect 295 6976 11944 6986
rect 12046 9686 12115 10493
rect 12149 10493 12151 10571
rect 12046 7712 12054 9686
rect 496 5313 1636 6976
rect 12046 6893 12115 7712
rect 2181 6751 7885 6752
rect 2134 6725 7885 6751
rect 2134 6668 2219 6725
rect 7862 6668 7885 6725
rect 2134 6593 7885 6668
rect 2134 6150 2288 6593
rect 7565 6151 7885 6593
rect 9855 6866 12115 6893
rect 9855 6841 10031 6866
rect 2134 5924 2503 6150
rect 2777 5924 3119 6150
rect 3393 5924 3735 6150
rect 4009 5924 4351 6150
rect 4625 5924 4967 6150
rect 5241 5924 5583 6150
rect 5857 5924 6199 6150
rect 6473 5924 6815 6150
rect 7565 6150 8009 6151
rect 7089 5924 8009 6150
rect 2134 5469 2288 5924
rect 7881 5469 8009 5924
rect 2134 5312 8009 5469
rect 2181 5311 8009 5312
rect 2181 5310 7900 5311
rect 7877 5206 8000 5207
rect 1020 5047 8000 5206
rect 1020 4611 1151 5047
rect 6591 4618 7453 5047
rect 1020 4449 1122 4611
rect 6591 4607 6796 4618
rect 1278 4605 6796 4607
rect 1278 4448 1661 4605
rect 1916 4448 2217 4605
rect 2472 4448 2773 4605
rect 3028 4448 3329 4605
rect 3584 4448 3885 4605
rect 4140 4448 4441 4605
rect 4696 4448 4997 4605
rect 5252 4448 5553 4605
rect 5808 4448 6109 4605
rect 6364 4449 6796 4605
rect 6952 4607 7453 4618
rect 7877 4607 8000 5047
rect 6952 4449 8000 4607
rect 6364 4448 8000 4449
rect 7877 4013 8000 4448
rect 127 199 210 4005
rect 1131 3963 8000 4013
rect 1131 3928 7905 3963
rect 1131 3873 1183 3928
rect 7858 3873 7905 3928
rect 9855 3943 9880 6841
rect 9945 6801 10031 6841
rect 11457 6817 12115 6866
rect 11457 6801 12149 6817
rect 9945 6777 12149 6801
rect 9945 6743 10048 6777
rect 12079 6743 12149 6777
rect 9945 6731 12149 6743
rect 9945 6695 10004 6731
rect 9945 4029 9963 6695
rect 9997 4029 10004 6695
rect 10519 6573 10924 6580
rect 10519 6444 10633 6573
rect 10519 5942 10924 6444
rect 11596 6250 12049 6252
rect 10193 5734 10924 5942
rect 11591 6249 12049 6250
rect 11591 6122 11623 6249
rect 11827 6122 12049 6249
rect 11591 6119 12049 6122
rect 11591 6023 11734 6119
rect 11591 5960 11616 6023
rect 11723 5960 11734 6023
rect 11591 5797 11734 5960
rect 11591 5767 12049 5797
rect 10452 5491 10924 5734
rect 11593 5722 12049 5767
rect 11593 5540 12049 5615
rect 10188 5476 10924 5491
rect 10188 5475 10813 5476
rect 10188 5248 10231 5475
rect 10404 5248 10813 5475
rect 11595 5396 11738 5540
rect 10188 5234 10813 5248
rect 11572 5388 11738 5396
rect 11572 5192 11601 5388
rect 11735 5192 11738 5388
rect 11572 5131 11738 5192
rect 11572 5057 12054 5131
rect 11576 5056 12054 5057
rect 11257 4826 11577 4957
rect 11624 4939 12054 5014
rect 10217 4685 10423 4687
rect 10217 4683 11590 4685
rect 11624 4683 11739 4939
rect 10217 4673 11739 4683
rect 10217 4513 10231 4673
rect 10408 4637 11739 4673
rect 10408 4513 12054 4637
rect 10217 4498 12054 4513
rect 9945 4017 10004 4029
rect 9945 3977 12149 4017
rect 9945 3943 10048 3977
rect 12078 3943 12149 3977
rect 9855 3909 12149 3943
rect 9855 3893 12115 3909
rect 1131 3854 7905 3873
rect 306 3771 11951 3789
rect 306 3768 5374 3771
rect 306 3689 1862 3768
rect 3521 3692 5374 3768
rect 7033 3692 11951 3771
rect 3521 3689 11951 3692
rect 306 3675 11951 3689
rect 306 3045 420 3675
rect 306 1084 319 3045
rect 413 1084 420 3045
rect 306 427 420 1084
rect 11837 3046 11951 3675
rect 11837 1085 11840 3046
rect 11934 1085 11951 3046
rect 11837 427 11951 1085
rect 306 313 11951 427
rect 12046 199 12115 3893
rect 127 153 12115 199
rect 86 127 12149 153
rect 86 93 153 127
rect 12089 93 12149 127
<< viali >>
rect 112 4005 127 7683
rect 127 4005 193 7683
rect 8302 6986 9743 7071
rect 12054 7712 12115 9686
rect 12115 7712 12142 9686
rect 2219 6668 7862 6725
rect 8319 6547 9723 6880
rect 2503 5924 2777 6151
rect 3119 5924 3393 6151
rect 3735 5924 4009 6151
rect 4351 5924 4625 6151
rect 4967 5924 5241 6151
rect 5583 5924 5857 6151
rect 6199 5924 6473 6151
rect 6815 5924 7089 6151
rect 1122 4442 1278 4611
rect 1661 4448 1916 4605
rect 2217 4448 2472 4605
rect 2773 4448 3028 4605
rect 3329 4448 3584 4605
rect 3885 4448 4140 4605
rect 4441 4448 4696 4605
rect 4997 4448 5252 4605
rect 5553 4448 5808 4605
rect 6109 4448 6364 4605
rect 6796 4449 6952 4618
rect 1183 3873 7858 3928
rect 8312 3923 9716 4256
rect 9880 3943 9945 6841
rect 10031 6801 11457 6866
rect 10633 6444 10929 6573
rect 11623 6122 11827 6249
rect 11616 5960 11723 6023
rect 10231 5248 10404 5475
rect 11601 5192 11735 5388
rect 10231 4513 10408 4673
rect 1862 3689 3521 3768
rect 5374 3692 7033 3771
rect 319 1084 413 3045
rect 11840 1085 11934 3046
<< metal1 >>
rect 514 9768 750 10200
rect 846 9768 1082 10200
rect 1178 9768 1414 10200
rect 1510 9768 1746 10200
rect 1842 9768 2078 10200
rect 2174 9768 2410 10200
rect 2506 9768 2742 10200
rect 2838 9768 3074 10200
rect 3170 9768 3406 10200
rect 3502 9768 3738 10200
rect 3834 9768 4070 10200
rect 4166 9768 4402 10200
rect 4498 9768 4734 10200
rect 4830 9768 5066 10200
rect 5162 9768 5398 10200
rect 5494 9768 5730 10200
rect 5826 9768 6062 10200
rect 6158 9768 6394 10200
rect 6490 9768 6726 10200
rect 6822 9768 7058 10200
rect 7154 9768 7390 10200
rect 7486 9768 7722 10200
rect 7818 9768 8054 10200
rect 8150 9768 8386 10200
rect 8482 9768 8718 10200
rect 8814 9768 9050 10200
rect 9146 9768 9382 10200
rect 9478 9768 9714 10200
rect 9810 9768 10046 10200
rect 10142 9768 10378 10200
rect 10474 9768 10710 10200
rect 10806 9768 11042 10200
rect 11138 9768 11374 10200
rect 11470 9768 11706 10200
rect 12048 9686 12148 9698
rect 12044 7712 12054 9686
rect 12142 7712 12152 9686
rect 12048 7700 12148 7712
rect 106 7683 199 7695
rect 102 4005 112 7683
rect 193 6463 203 7683
rect 513 6641 588 7601
rect 680 7168 916 7600
rect 1012 7168 1248 7600
rect 1344 7168 1580 7600
rect 1676 7168 1912 7600
rect 2008 7168 2244 7600
rect 2340 7168 2576 7600
rect 2672 7168 2908 7600
rect 3004 7168 3240 7600
rect 3336 7168 3572 7600
rect 3668 7168 3904 7600
rect 4000 7168 4236 7600
rect 4332 7168 4568 7600
rect 4664 7168 4900 7600
rect 4996 7168 5232 7600
rect 5328 7168 5564 7600
rect 5660 7168 5896 7600
rect 5992 7168 6228 7600
rect 6324 7168 6560 7600
rect 6656 7168 6892 7600
rect 6988 7168 7224 7600
rect 7320 7168 7556 7600
rect 7652 7168 7888 7600
rect 7984 7168 8220 7600
rect 8316 7168 8552 7600
rect 8648 7168 8884 7600
rect 8980 7168 9216 7600
rect 9312 7168 9548 7600
rect 9644 7168 9880 7600
rect 9976 7168 10212 7600
rect 10308 7168 10544 7600
rect 10640 7168 10876 7600
rect 10972 7168 11208 7600
rect 11304 7168 11540 7600
rect 627 7080 1828 7083
rect 8285 7080 9768 7090
rect 627 7071 9768 7080
rect 627 7069 8302 7071
rect 627 6942 654 7069
rect 1795 6986 8302 7069
rect 9743 6986 9768 7071
rect 1795 6942 9768 6986
rect 627 6925 9768 6942
rect 807 6924 9768 6925
rect 8285 6901 9768 6924
rect 9837 6999 11494 7024
rect 9837 6901 9877 6999
rect 11458 6901 11494 6999
rect 8285 6880 9767 6901
rect 2137 6818 7913 6848
rect 2137 6753 2190 6818
rect 7886 6753 7913 6818
rect 2137 6725 7913 6753
rect 2137 6668 2219 6725
rect 7862 6668 7913 6725
rect 2137 6658 7913 6668
rect 513 6590 1839 6641
rect 193 5310 1632 6463
rect 193 4005 203 5310
rect 1439 4946 1449 4967
rect 1194 4623 1278 4871
rect 1348 4720 1376 4937
rect 1384 4906 1449 4946
rect 1439 4905 1449 4906
rect 1606 4905 1616 4967
rect 1116 4611 1284 4623
rect 1112 4442 1122 4611
rect 1278 4442 1288 4611
rect 1116 4430 1284 4442
rect 1454 4129 1486 4868
rect 1788 4790 1839 6590
rect 8285 6547 8319 6880
rect 9723 6547 9767 6880
rect 2373 6475 6862 6522
rect 8285 6506 9767 6547
rect 9837 6866 11494 6901
rect 9837 6841 10031 6866
rect 2373 5696 2420 6475
rect 2483 6265 2514 6475
rect 2573 6157 2673 6415
rect 2491 6151 2789 6157
rect 2491 5924 2503 6151
rect 2777 5924 2789 6151
rect 2491 5918 2789 5924
rect 2336 5649 2420 5696
rect 1960 5063 1970 5084
rect 1903 5022 1970 5063
rect 2127 5063 2137 5084
rect 2127 5026 2217 5063
rect 2127 5022 2137 5026
rect 1903 4722 1940 5022
rect 1649 4605 1928 4611
rect 1649 4448 1661 4605
rect 1916 4448 1928 4605
rect 1649 4442 1928 4448
rect 1747 4185 1831 4442
rect 1904 4129 1937 4328
rect 2009 4129 2049 4879
rect 2180 4752 2217 5026
rect 2336 4786 2383 5649
rect 2482 5088 2514 5802
rect 2588 5652 2692 5918
rect 2985 5653 3029 6422
rect 3099 6265 3130 6475
rect 3189 6157 3289 6415
rect 3107 6151 3405 6157
rect 3107 5924 3119 6151
rect 3393 5924 3405 6151
rect 3107 5918 3405 5924
rect 3092 5328 3131 5807
rect 2993 5163 3003 5328
rect 3060 5286 3131 5328
rect 3190 5516 3229 5734
rect 3601 5653 3645 6422
rect 3715 6265 3746 6475
rect 3805 6157 3905 6415
rect 3723 6151 4021 6157
rect 3723 5924 3735 6151
rect 4009 5924 4021 6151
rect 3723 5918 4021 5924
rect 3190 5426 3204 5516
rect 3414 5426 3424 5516
rect 3190 5326 3229 5426
rect 3708 5326 3747 5807
rect 3190 5287 3747 5326
rect 3819 5516 3858 5738
rect 4217 5653 4261 6422
rect 4331 6265 4362 6475
rect 4421 6157 4521 6415
rect 4339 6151 4637 6157
rect 4339 5924 4351 6151
rect 4625 5924 4637 6151
rect 4339 5918 4637 5924
rect 3819 5426 3835 5516
rect 4045 5426 4055 5516
rect 3819 5328 3858 5426
rect 4324 5328 4363 5807
rect 3819 5289 4363 5328
rect 4445 5516 4484 5745
rect 4833 5653 4877 6422
rect 4947 6265 4978 6475
rect 5037 6157 5137 6415
rect 4955 6151 5253 6157
rect 4955 5924 4967 6151
rect 5241 5924 5253 6151
rect 4955 5918 5253 5924
rect 4445 5426 4467 5516
rect 4677 5426 4687 5516
rect 4445 5328 4484 5426
rect 4940 5328 4979 5807
rect 4445 5289 4979 5328
rect 5048 5516 5087 5737
rect 5449 5653 5493 6422
rect 5563 6265 5594 6475
rect 5653 6157 5753 6415
rect 5571 6151 5869 6157
rect 5571 5924 5583 6151
rect 5857 5924 5869 6151
rect 5571 5918 5869 5924
rect 5048 5426 5071 5516
rect 5281 5426 5291 5516
rect 5048 5328 5087 5426
rect 5556 5328 5595 5807
rect 5048 5289 5595 5328
rect 5672 5498 5711 5744
rect 6065 5653 6109 6422
rect 6179 6265 6210 6475
rect 6269 6157 6369 6415
rect 6187 6151 6485 6157
rect 6187 5924 6199 6151
rect 6473 5924 6485 6151
rect 6187 5918 6485 5924
rect 5874 5498 5884 5516
rect 5672 5442 5884 5498
rect 5672 5328 5711 5442
rect 5874 5426 5884 5442
rect 6094 5426 6104 5516
rect 6172 5328 6211 5807
rect 5672 5289 6211 5328
rect 6283 5328 6322 5741
rect 6681 5653 6725 6422
rect 6795 6265 6826 6475
rect 6885 6157 6985 6415
rect 7502 6173 7512 6272
rect 7872 6173 7882 6272
rect 6803 6151 7101 6157
rect 6803 5924 6815 6151
rect 7089 5924 7101 6151
rect 6803 5918 7101 5924
rect 6788 5328 6827 5807
rect 6905 5332 6944 5744
rect 7511 5666 7595 6173
rect 8020 5967 8030 5988
rect 7758 5929 8030 5967
rect 7656 5513 7700 5824
rect 7203 5469 7700 5513
rect 6283 5289 6827 5328
rect 3060 5163 3070 5286
rect 2472 5026 2482 5088
rect 2639 5026 2649 5088
rect 2459 4752 2496 4959
rect 2180 4715 2496 4752
rect 2205 4605 2484 4611
rect 2205 4448 2217 4605
rect 2472 4448 2484 4605
rect 2205 4442 2484 4448
rect 2303 4431 2395 4442
rect 2311 4188 2395 4431
rect 2461 4130 2494 4333
rect 2561 4188 2603 4877
rect 2904 4681 2946 4874
rect 3016 4720 3055 5163
rect 3190 5015 3229 5287
rect 3128 4976 3229 5015
rect 3128 4787 3167 4976
rect 3460 4681 3502 4874
rect 3572 4720 3611 5287
rect 3819 5016 3858 5289
rect 3679 4977 3858 5016
rect 3679 4781 3718 4977
rect 4016 4681 4058 4874
rect 4128 4720 4167 5289
rect 4445 5018 4484 5289
rect 4235 4979 4484 5018
rect 4235 4789 4274 4979
rect 4572 4681 4614 4874
rect 4684 4720 4723 5289
rect 5048 5021 5087 5289
rect 4789 4982 5087 5021
rect 4789 4781 4828 4982
rect 5128 4681 5170 4874
rect 5240 4720 5279 5289
rect 5672 5020 5711 5289
rect 5347 4981 5711 5020
rect 5347 4782 5386 4981
rect 5684 4681 5726 4874
rect 5796 4720 5835 5289
rect 6283 5027 6322 5289
rect 5910 4988 6322 5027
rect 5910 4786 5949 4988
rect 6240 4681 6282 4874
rect 6352 4720 6391 5289
rect 6892 5167 6902 5332
rect 6959 5290 6969 5332
rect 7203 5290 7247 5469
rect 6959 5223 7247 5290
rect 6959 5167 6969 5223
rect 6905 5032 6944 5167
rect 6457 4993 6944 5032
rect 6457 4787 6496 4993
rect 2904 4639 3159 4681
rect 3460 4639 3715 4681
rect 4016 4639 4271 4681
rect 4572 4639 4827 4681
rect 5128 4639 5383 4681
rect 5684 4639 5939 4681
rect 6240 4639 6495 4681
rect 2761 4605 3040 4611
rect 2761 4448 2773 4605
rect 3028 4448 3040 4605
rect 2761 4442 3040 4448
rect 2859 4431 2951 4442
rect 2867 4188 2951 4431
rect 3017 4130 3050 4333
rect 3117 4188 3159 4639
rect 3317 4605 3596 4611
rect 3317 4448 3329 4605
rect 3584 4448 3596 4605
rect 3317 4442 3596 4448
rect 3415 4431 3507 4442
rect 3423 4188 3507 4431
rect 3573 4130 3606 4333
rect 3673 4188 3715 4639
rect 3873 4605 4152 4611
rect 3873 4448 3885 4605
rect 4140 4448 4152 4605
rect 3873 4442 4152 4448
rect 3971 4431 4063 4442
rect 3979 4188 4063 4431
rect 4129 4130 4162 4333
rect 4229 4188 4271 4639
rect 4429 4605 4708 4611
rect 4429 4448 4441 4605
rect 4696 4448 4708 4605
rect 4429 4442 4708 4448
rect 4527 4431 4619 4442
rect 4535 4188 4619 4431
rect 4685 4130 4718 4333
rect 4785 4188 4827 4639
rect 4985 4605 5264 4611
rect 4985 4448 4997 4605
rect 5252 4448 5264 4605
rect 4985 4442 5264 4448
rect 5083 4431 5175 4442
rect 5091 4188 5175 4431
rect 5241 4130 5274 4333
rect 5341 4188 5383 4639
rect 5541 4605 5820 4611
rect 5541 4448 5553 4605
rect 5808 4448 5820 4605
rect 5541 4442 5820 4448
rect 5639 4431 5731 4442
rect 5647 4188 5731 4431
rect 5797 4130 5830 4333
rect 5897 4188 5939 4639
rect 6097 4605 6376 4611
rect 6097 4448 6109 4605
rect 6364 4448 6376 4605
rect 6097 4442 6376 4448
rect 6195 4431 6287 4442
rect 6203 4188 6287 4431
rect 6353 4130 6386 4333
rect 6453 4188 6495 4639
rect 6790 4618 6958 4630
rect 6790 4613 6796 4618
rect 6656 4605 6796 4613
rect 6656 4448 6665 4605
rect 6952 4449 6958 4618
rect 6920 4448 6958 4449
rect 6656 4439 6958 4448
rect 6790 4437 6958 4439
rect 7203 4447 7247 5223
rect 7544 4623 7582 4860
rect 7649 4743 7685 4933
rect 7758 4785 7796 5929
rect 8020 5910 8030 5929
rect 8221 5910 8231 5988
rect 8050 5145 8329 5179
rect 8050 4961 8084 5145
rect 7930 4897 7940 4961
rect 8127 4897 8137 4961
rect 7649 4707 8069 4743
rect 8033 4638 8069 4707
rect 7544 4585 7795 4623
rect 8033 4599 8097 4638
rect 6824 4274 6908 4437
rect 7203 4404 7690 4447
rect 7261 4403 7690 4404
rect 6824 4273 7584 4274
rect 6824 4191 7594 4273
rect 6824 4190 7482 4191
rect 1454 4081 6404 4129
rect 7646 4124 7690 4403
rect 7757 4190 7795 4585
rect 8087 4574 8097 4599
rect 8284 4574 8294 4638
rect 9837 4316 9880 6841
rect 9725 4306 9880 4316
rect 8268 4256 9880 4306
rect 106 3993 199 4005
rect 1129 3928 7903 4013
rect 1129 3873 1183 3928
rect 7858 3873 7903 3928
rect 8268 3923 8312 4256
rect 9716 3943 9880 4256
rect 9945 6801 10031 6841
rect 11457 6801 11494 6866
rect 9945 6774 11494 6801
rect 9945 3943 10014 6774
rect 11658 6702 11733 7607
rect 10494 6627 11733 6702
rect 10267 6483 10277 6555
rect 10453 6483 10463 6555
rect 10254 5988 10307 6188
rect 10391 6102 10453 6483
rect 10065 5916 10075 5988
rect 10251 5934 10307 5988
rect 10251 5916 10261 5934
rect 10352 5780 10384 6064
rect 10240 5708 10250 5780
rect 10426 5708 10436 5780
rect 10352 5641 10384 5643
rect 10212 5569 10222 5641
rect 10398 5569 10408 5641
rect 10217 5475 10423 5493
rect 10217 5248 10231 5475
rect 10404 5248 10423 5475
rect 10217 4673 10423 5248
rect 10217 4513 10231 4673
rect 10408 4513 10423 4673
rect 10217 4500 10423 4513
rect 10494 4131 10569 6627
rect 10621 6573 10941 6579
rect 10621 6444 10633 6573
rect 10929 6444 10941 6573
rect 11864 6564 12242 7121
rect 10621 6438 10941 6444
rect 11142 6554 12242 6564
rect 11142 6455 11153 6554
rect 11513 6455 12242 6554
rect 11142 6364 12242 6455
rect 10638 6177 10648 6276
rect 11008 6177 11018 6276
rect 11142 6249 11839 6364
rect 10644 4934 10806 6177
rect 11142 6122 11623 6249
rect 11827 6122 11839 6249
rect 11142 6116 11839 6122
rect 11142 6039 11629 6116
rect 11142 6023 11838 6039
rect 11142 5960 11616 6023
rect 11723 5960 11838 6023
rect 11142 5945 11838 5960
rect 11142 5943 11342 5945
rect 11829 5944 11838 5945
rect 11938 5938 11986 6044
rect 11938 5890 12060 5938
rect 11818 5829 11904 5883
rect 11489 5655 11499 5672
rect 11428 5600 11499 5655
rect 11675 5663 11685 5672
rect 11818 5663 11859 5829
rect 11675 5614 11859 5663
rect 11675 5600 11685 5614
rect 11428 5290 11466 5600
rect 11818 5431 11859 5614
rect 11887 5613 11897 5782
rect 11966 5613 11976 5782
rect 11910 5530 11976 5613
rect 11595 5388 11741 5400
rect 11338 5252 11466 5290
rect 11338 5136 11376 5252
rect 11503 5222 11601 5388
rect 11435 5192 11601 5222
rect 11735 5192 11841 5388
rect 11435 5190 11841 5192
rect 11435 5180 11741 5190
rect 11435 5140 11715 5180
rect 11253 5026 11263 5098
rect 11439 5026 11449 5098
rect 11503 4934 11715 5140
rect 11935 5127 11976 5530
rect 10644 4734 11715 4934
rect 11787 5086 11976 5127
rect 11787 4786 11828 5086
rect 12012 5038 12060 5890
rect 11939 4990 12060 5038
rect 11939 4786 11987 4990
rect 11155 4391 11715 4734
rect 11777 4671 11787 4730
rect 11973 4671 11983 4730
rect 11155 4191 12242 4391
rect 10494 4056 11733 4131
rect 9716 3923 10014 3943
rect 8268 3892 10014 3923
rect 1129 3856 7903 3873
rect 1850 3768 3533 3774
rect 1850 3689 1862 3768
rect 3521 3689 3533 3768
rect 1850 3683 3533 3689
rect 5362 3771 7045 3777
rect 5362 3692 5374 3771
rect 7033 3692 7045 3771
rect 5362 3686 7045 3692
rect 86 3543 605 3550
rect 86 3134 100 3543
rect 351 3134 605 3543
rect 86 3118 605 3134
rect 700 3118 936 3550
rect 1032 3118 1268 3550
rect 1364 3118 1600 3550
rect 1696 3118 1932 3550
rect 2028 3118 2264 3550
rect 2360 3118 2596 3550
rect 2692 3118 2928 3550
rect 3024 3118 3260 3550
rect 3356 3118 3592 3550
rect 3688 3118 3924 3550
rect 4020 3118 4256 3550
rect 4352 3118 4588 3550
rect 4684 3118 4920 3550
rect 5016 3118 5252 3550
rect 5348 3118 5584 3550
rect 5680 3118 5916 3550
rect 6012 3118 6248 3550
rect 6344 3118 6580 3550
rect 6676 3118 6912 3550
rect 7008 3118 7244 3550
rect 7340 3118 7576 3550
rect 7672 3118 7908 3550
rect 8004 3118 8240 3550
rect 8336 3118 8572 3550
rect 8668 3118 8904 3550
rect 9000 3118 9236 3550
rect 9332 3118 9568 3550
rect 9664 3118 9900 3550
rect 9996 3118 10232 3550
rect 10328 3118 10564 3550
rect 10660 3118 10896 3550
rect 10992 3118 11228 3550
rect 11324 3118 11560 3550
rect 11658 3115 11733 4056
rect 11864 3634 12242 4191
rect 313 3045 419 3057
rect 11834 3046 11940 3058
rect 309 1084 319 3045
rect 413 1084 423 3045
rect 11830 1085 11840 3046
rect 11934 1085 11944 3046
rect 313 1072 419 1084
rect 11834 1073 11940 1085
rect 534 518 770 950
rect 866 518 1102 950
rect 1198 518 1434 950
rect 1530 518 1766 950
rect 1862 518 2098 950
rect 2194 518 2430 950
rect 2526 518 2762 950
rect 2858 518 3094 950
rect 3190 518 3426 950
rect 3522 518 3758 950
rect 3854 518 4090 950
rect 4186 518 4422 950
rect 4518 518 4754 950
rect 4850 518 5086 950
rect 5182 518 5418 950
rect 5514 518 5750 950
rect 5846 518 6082 950
rect 6178 518 6414 950
rect 6510 518 6746 950
rect 6842 518 7078 950
rect 7174 518 7410 950
rect 7506 518 7742 950
rect 7838 518 8074 950
rect 8170 518 8406 950
rect 8502 518 8738 950
rect 8834 518 9070 950
rect 9166 518 9402 950
rect 9498 518 9734 950
rect 9830 518 10066 950
rect 10162 518 10398 950
rect 10494 518 10730 950
rect 10826 518 11062 950
rect 11158 518 11394 950
rect 11490 518 11726 950
<< via1 >>
rect 12054 7712 12142 9686
rect 112 4005 193 7683
rect 654 6942 1795 7069
rect 9877 6901 11458 6999
rect 2190 6753 7886 6818
rect 1449 4905 1606 4967
rect 1122 4442 1278 4611
rect 8319 6547 9723 6880
rect 2503 5924 2777 6151
rect 1970 5022 2127 5084
rect 1661 4448 1916 4605
rect 3119 5924 3393 6151
rect 3003 5163 3060 5328
rect 3735 5924 4009 6151
rect 3204 5426 3414 5516
rect 4351 5924 4625 6151
rect 3835 5426 4045 5516
rect 4967 5924 5241 6151
rect 4467 5426 4677 5516
rect 5583 5924 5857 6151
rect 5071 5426 5281 5516
rect 6199 5924 6473 6151
rect 5884 5426 6094 5516
rect 7512 6173 7872 6272
rect 6815 5924 7089 6151
rect 2482 5026 2639 5088
rect 2217 4448 2472 4605
rect 6902 5167 6959 5332
rect 2773 4448 3028 4605
rect 3329 4448 3584 4605
rect 3885 4448 4140 4605
rect 4441 4448 4696 4605
rect 4997 4448 5252 4605
rect 5553 4448 5808 4605
rect 6109 4448 6364 4605
rect 6665 4449 6796 4605
rect 6796 4449 6920 4605
rect 6665 4448 6920 4449
rect 8030 5910 8221 5988
rect 7940 4897 8127 4961
rect 8097 4574 8284 4638
rect 1183 3873 7858 3928
rect 8312 3923 9716 4256
rect 10277 6483 10453 6555
rect 10075 5916 10251 5988
rect 10250 5708 10426 5780
rect 10222 5569 10398 5641
rect 10633 6444 10929 6573
rect 11153 6455 11513 6554
rect 10648 6177 11008 6276
rect 11499 5600 11675 5672
rect 11897 5613 11966 5782
rect 11263 5026 11439 5098
rect 11787 4671 11973 4730
rect 1862 3689 3521 3768
rect 5374 3692 7033 3771
rect 100 3134 351 3543
rect 319 1084 413 3045
rect 11840 1085 11934 3046
<< metal2 >>
rect 12054 9695 12142 9696
rect 0 9686 12242 9695
rect 0 7712 12054 9686
rect 12142 7712 12242 9686
rect 0 7701 12242 7712
rect 92 7683 358 7701
rect 92 4005 112 7683
rect 193 4005 358 7683
rect 627 7069 1828 7083
rect 627 7065 654 7069
rect 92 3543 358 4005
rect 92 3134 100 3543
rect 351 3134 358 3543
rect 92 3128 358 3134
rect 625 6942 654 7065
rect 1795 6942 1828 7069
rect 625 6925 1828 6942
rect 625 6464 1175 6925
rect 2453 6865 4111 7701
rect 5409 6865 7067 7701
rect 8285 6901 9768 7090
rect 9837 6999 11494 7701
rect 9837 6901 9877 6999
rect 11458 6901 11494 6999
rect 8285 6880 9767 6901
rect 9837 6882 11494 6901
rect 2119 6818 7954 6865
rect 2119 6753 2190 6818
rect 7886 6753 7954 6818
rect 2119 6655 7954 6753
rect 625 5307 1635 6464
rect 2453 6199 4111 6655
rect 5409 6199 7067 6655
rect 8285 6547 8319 6880
rect 9723 6547 9767 6880
rect 10633 6574 10929 6583
rect 8285 6506 9767 6547
rect 10263 6573 11518 6574
rect 10263 6555 10633 6573
rect 10263 6483 10277 6555
rect 10453 6483 10633 6555
rect 10263 6444 10633 6483
rect 10929 6554 11518 6573
rect 10929 6455 11153 6554
rect 11513 6455 11518 6554
rect 10929 6444 11518 6455
rect 10263 6442 11518 6444
rect 10633 6434 10929 6442
rect 7512 6274 7872 6282
rect 10648 6276 11008 6286
rect 7512 6272 10648 6274
rect 2131 6151 7166 6199
rect 7872 6177 10648 6272
rect 7872 6176 11008 6177
rect 7512 6163 7872 6173
rect 10648 6167 11008 6176
rect 2131 5924 2503 6151
rect 2777 5924 3119 6151
rect 3393 5924 3735 6151
rect 4009 5924 4351 6151
rect 4625 5924 4967 6151
rect 5241 5924 5583 6151
rect 5857 5924 6199 6151
rect 6473 5924 6815 6151
rect 7089 5924 7166 6151
rect 2131 5883 7166 5924
rect 8030 5988 8221 5998
rect 10075 5988 10251 5998
rect 8221 5929 9972 5973
rect 10074 5929 10075 5973
rect 8030 5900 8221 5910
rect 9928 5876 9972 5929
rect 10251 5929 11574 5973
rect 10075 5906 10251 5916
rect 9928 5832 11424 5876
rect 10250 5780 10426 5790
rect 10250 5698 10426 5708
rect 11380 5654 11424 5832
rect 11530 5759 11574 5929
rect 11897 5782 11966 5792
rect 11530 5715 11897 5759
rect 11499 5672 11675 5682
rect 10222 5641 10398 5651
rect 2521 5592 2619 5602
rect 3587 5592 3685 5602
rect 3204 5523 3414 5526
rect 2619 5516 3414 5523
rect 2619 5426 3204 5516
rect 2619 5418 3414 5426
rect 3204 5416 3414 5418
rect 2521 5367 2619 5377
rect 4653 5592 4751 5602
rect 3685 5526 3851 5527
rect 3685 5516 4045 5526
rect 3685 5426 3835 5516
rect 3685 5417 4045 5426
rect 3835 5416 4045 5417
rect 4467 5516 4653 5526
rect 5719 5592 5817 5602
rect 4467 5416 4653 5426
rect 3587 5367 3685 5377
rect 5071 5516 5719 5526
rect 5281 5426 5719 5516
rect 5071 5417 5719 5426
rect 5071 5416 5281 5417
rect 4653 5367 4751 5377
rect 6785 5592 6883 5602
rect 6082 5526 6785 5527
rect 5884 5516 6785 5526
rect 6094 5426 6785 5516
rect 5884 5417 6785 5426
rect 5884 5416 6094 5417
rect 5719 5367 5817 5377
rect 6785 5367 6883 5377
rect 3003 5328 3060 5338
rect 625 4644 1175 5307
rect 6902 5332 6959 5342
rect 3060 5220 6902 5261
rect 3003 5153 3060 5163
rect 6902 5157 6959 5167
rect 1970 5084 2127 5094
rect 2482 5088 2639 5098
rect 1932 5023 1970 5084
rect 2127 5026 2482 5084
rect 2639 5026 8263 5084
rect 2127 5023 8263 5026
rect 1970 5012 2127 5022
rect 2482 5016 2639 5023
rect 1449 4967 1606 4977
rect 7930 4961 8127 4971
rect 7930 4950 7940 4961
rect 1606 4905 7940 4950
rect 1449 4895 1606 4905
rect 7940 4887 8127 4897
rect 8202 4926 8263 5023
rect 8202 4865 8538 4926
rect 625 4611 7135 4644
rect 8097 4639 8284 4648
rect 9688 4639 9753 5600
rect 11380 5610 11499 5654
rect 12042 5759 12242 5830
rect 11966 5715 12242 5759
rect 12042 5630 12242 5715
rect 11897 5603 11966 5613
rect 11499 5590 11675 5600
rect 10222 5559 10398 5569
rect 11016 5391 11569 5445
rect 11263 5098 11439 5108
rect 11515 5086 11569 5391
rect 11439 5039 11569 5086
rect 11263 5016 11439 5026
rect 11515 4913 11569 5039
rect 12042 4913 12242 4986
rect 11515 4859 12242 4913
rect 11854 4740 11910 4859
rect 12042 4786 12242 4859
rect 11787 4730 11973 4740
rect 11787 4661 11973 4671
rect 625 4442 1122 4611
rect 1278 4605 7135 4611
rect 1278 4448 1661 4605
rect 1916 4448 2217 4605
rect 2472 4448 2773 4605
rect 3028 4448 3329 4605
rect 3584 4448 3885 4605
rect 4140 4448 4441 4605
rect 4696 4448 4997 4605
rect 5252 4448 5553 4605
rect 5808 4448 6109 4605
rect 6364 4448 6665 4605
rect 6920 4448 7135 4605
rect 8095 4638 9753 4639
rect 8095 4574 8097 4638
rect 8284 4574 9753 4638
rect 8097 4564 8284 4574
rect 1278 4442 7135 4448
rect 625 4342 7135 4442
rect 625 4038 1175 4342
rect 1861 4038 3520 4342
rect 5375 4038 7034 4342
rect 8268 4256 9750 4306
rect 625 3928 7930 4038
rect 625 3873 1183 3928
rect 7858 3873 7930 3928
rect 8268 3923 8312 4256
rect 9716 3923 9750 4256
rect 8268 3892 9750 3923
rect 625 3824 7930 3873
rect 625 3062 1175 3824
rect 1861 3768 3521 3824
rect 1861 3689 1862 3768
rect 1861 3679 3521 3689
rect 5374 3771 7034 3824
rect 7033 3692 7034 3771
rect 5374 3682 7034 3692
rect 1861 3062 3520 3679
rect 5375 3062 7034 3682
rect 0 3046 12242 3062
rect 0 3045 11840 3046
rect 0 1084 319 3045
rect 413 3008 11840 3045
rect 413 2741 3091 3008
rect 7477 2741 11840 3008
rect 413 1085 11840 2741
rect 11934 1085 12242 3046
rect 413 1084 12242 1085
rect 0 1068 12242 1084
<< via2 >>
rect 2521 5377 2619 5592
rect 3587 5377 3685 5592
rect 4653 5516 4751 5592
rect 4653 5426 4677 5516
rect 4677 5426 4751 5516
rect 4653 5377 4751 5426
rect 5719 5377 5817 5592
rect 6785 5377 6883 5592
rect 3091 2741 7477 3008
<< metal3 >>
rect 2511 5592 2629 5597
rect 2511 5377 2521 5592
rect 2619 5377 2629 5592
rect 2511 5372 2629 5377
rect 3577 5592 3695 5597
rect 3577 5377 3587 5592
rect 3685 5377 3695 5592
rect 3577 5372 3695 5377
rect 4643 5592 4761 5597
rect 4643 5377 4653 5592
rect 4751 5377 4761 5592
rect 4643 5372 4761 5377
rect 5709 5592 5827 5597
rect 5709 5377 5719 5592
rect 5817 5377 5827 5592
rect 5709 5372 5827 5377
rect 6775 5592 6893 5597
rect 6775 5377 6785 5592
rect 6883 5377 6893 5592
rect 6775 5372 6893 5377
rect 3204 3930 3298 5210
rect 4270 3930 4364 5210
rect 5336 3931 5430 5211
rect 6402 3931 6496 5211
rect 3094 3571 3104 3821
rect 3202 3571 3212 3821
rect 3094 3013 3212 3571
rect 4160 3571 4170 3821
rect 4268 3571 4278 3821
rect 4160 3013 4278 3571
rect 5226 3571 5236 3821
rect 5334 3571 5344 3821
rect 5226 3013 5344 3571
rect 6292 3571 6302 3821
rect 6400 3571 6410 3821
rect 6292 3013 6410 3571
rect 7358 3571 7368 3821
rect 7466 3571 7476 3821
rect 7358 3013 7476 3571
rect 3081 3008 7487 3013
rect 3081 2741 3091 3008
rect 7477 2741 7487 3008
rect 3081 2736 7487 2741
<< via3 >>
rect 2521 5377 2619 5592
rect 3587 5377 3685 5592
rect 4653 5377 4751 5592
rect 5719 5377 5817 5592
rect 6785 5377 6883 5592
rect 3104 3571 3202 3821
rect 4170 3571 4268 3821
rect 5236 3571 5334 3821
rect 6302 3571 6400 3821
rect 7368 3571 7466 3821
<< metal4 >>
rect 2510 5592 2630 5598
rect 2510 5377 2521 5592
rect 2619 5377 2630 5592
rect 2510 5370 2630 5377
rect 3576 5592 3696 5598
rect 3576 5377 3587 5592
rect 3685 5377 3696 5592
rect 3576 5370 3696 5377
rect 4642 5592 4762 5598
rect 4642 5377 4653 5592
rect 4751 5377 4762 5592
rect 4642 5370 4762 5377
rect 5708 5592 5828 5598
rect 5708 5377 5719 5592
rect 5817 5377 5828 5592
rect 5708 5370 5828 5377
rect 6774 5592 6894 5598
rect 6774 5377 6785 5592
rect 6883 5377 6894 5592
rect 6774 5370 6894 5377
rect 2521 4328 2619 5370
rect 3587 4328 3685 5370
rect 4653 4328 4751 5370
rect 5719 4328 5817 5370
rect 6785 4328 6883 5370
rect 3104 3822 3202 4080
rect 4170 3822 4268 4080
rect 5236 3822 5334 4080
rect 6302 3822 6400 4080
rect 7368 3822 7466 4080
rect 3103 3821 3203 3822
rect 3103 3571 3104 3821
rect 3202 3571 3203 3821
rect 3103 3570 3203 3571
rect 4169 3821 4269 3822
rect 4169 3571 4170 3821
rect 4268 3571 4269 3821
rect 4169 3570 4269 3571
rect 5235 3821 5335 3822
rect 5235 3571 5236 3821
rect 5334 3571 5335 3821
rect 5235 3570 5335 3571
rect 6301 3821 6401 3822
rect 6301 3571 6302 3821
rect 6400 3571 6401 3821
rect 6301 3570 6401 3571
rect 7367 3821 7467 3822
rect 7367 3571 7368 3821
rect 7466 3571 7467 3821
rect 7367 3570 7467 3571
use sky130_fd_pr__diode_pw2nd_05v5_FT76RJ  D3
timestamp 1699295625
transform 1 0 10339 0 1 5604
box -183 -183 183 183
use level_shifter  level_shifter_0
timestamp 1699295625
transform -1 0 10932 0 -1 4214
box -422 -2544 2736 144
use sky130_fd_pr__cap_mim_m3_1_AZFCP3  sky130_fd_pr__cap_mim_m3_1_AZFCP3_1
timestamp 1699295625
transform 1 0 6982 0 1 4571
box -486 -640 486 640
use sky130_fd_pr__nfet_01v8_L9WNCD  sky130_fd_pr__nfet_01v8_L9WNCD_0
timestamp 1699295625
transform 1 0 11875 0 1 5958
box -211 -229 211 229
use sky130_fd_pr__pfet_01v8_2Z69BZ  sky130_fd_pr__pfet_01v8_2Z69BZ_0
timestamp 1699295625
transform 1 0 11402 0 1 5145
box -211 -226 211 226
use sky130_fd_pr__pfet_01v8_LGS3BL  sky130_fd_pr__pfet_01v8_LGS3BL_0
timestamp 1699295625
transform 1 0 11878 0 -1 5325
box -211 -284 211 284
use sky130_fd_pr__res_xhigh_po_0p35_DEAPHQ  sky130_fd_pr__res_xhigh_po_0p35_DEAPHQ_0
timestamp 1699295625
transform 1 0 6130 0 1 2034
box -5762 -1682 5762 1682
use sky130_fd_pr__res_xhigh_po_0p35_DEAPHQ  sky130_fd_pr__res_xhigh_po_0p35_DEAPHQ_1
timestamp 1699295625
transform 1 0 6110 0 1 8684
box -5762 -1682 5762 1682
use sky130_fd_pr__cap_mim_m3_1_AZFCP3  XC1
timestamp 1699295625
transform 1 0 2718 0 1 4570
box -486 -640 486 640
use sky130_fd_pr__cap_mim_m3_1_AZFCP3  XC2
timestamp 1699295625
transform 1 0 3784 0 1 4570
box -486 -640 486 640
use sky130_fd_pr__cap_mim_m3_1_AZFCP3  XC3
timestamp 1699295625
transform 1 0 4850 0 1 4571
box -486 -640 486 640
use sky130_fd_pr__cap_mim_m3_1_AZFCP3  XC4
timestamp 1699295625
transform 1 0 5916 0 1 4571
box -486 -640 486 640
use sky130_fd_pr__nfet_g5v0d10v5_6XHUDR  XM1
timestamp 1699295625
transform 1 0 3032 0 1 4830
box -278 -300 278 300
use sky130_fd_pr__pfet_g5v0d10v5_6ELFTH  XM2
timestamp 1699295625
transform 1 0 3114 0 1 5695
box -308 -339 308 339
use sky130_fd_pr__pfet_g5v0d10v5_6ELFTH  XM3
timestamp 1699295625
transform 1 0 3730 0 1 5695
box -308 -339 308 339
use sky130_fd_pr__nfet_g5v0d10v5_6XHUDR  XM4
timestamp 1699295625
transform 1 0 3588 0 1 4830
box -278 -300 278 300
use sky130_fd_pr__nfet_01v8_L9WNCD  XM5
timestamp 1699295625
transform 1 0 11882 0 1 4794
box -211 -229 211 229
use sky130_fd_pr__pfet_g5v0d10v5_6ELFTH  XM7
timestamp 1699295625
transform 1 0 4962 0 1 5695
box -308 -339 308 339
use sky130_fd_pr__nfet_g5v0d10v5_6XHUDR  XM8
timestamp 1699295625
transform 1 0 4700 0 1 4830
box -278 -300 278 300
use sky130_fd_pr__pfet_g5v0d10v5_6ELFTH  XM9
timestamp 1699295625
transform 1 0 4346 0 1 5695
box -308 -339 308 339
use sky130_fd_pr__nfet_g5v0d10v5_6XHUDR  XM10
timestamp 1699295625
transform 1 0 4144 0 1 4830
box -278 -300 278 300
use sky130_fd_pr__pfet_g5v0d10v5_6ELFTH  XM11
timestamp 1699295625
transform 1 0 7680 0 1 5695
box -308 -339 308 339
use sky130_fd_pr__nfet_g5v0d10v5_6XHUDR  XM12
timestamp 1699295625
transform 1 0 7668 0 1 4228
box -278 -300 278 300
use sky130_fd_pr__nfet_g5v0d10v5_6XHUDR  XM13
timestamp 1699295625
transform 1 0 7668 0 1 4828
box -278 -300 278 300
use sky130_fd_pr__pfet_g5v0d10v5_6ELFTH  XM15
timestamp 1699295625
transform 1 0 5578 0 1 5695
box -308 -339 308 339
use sky130_fd_pr__nfet_g5v0d10v5_6XHUDR  XM16
timestamp 1699295625
transform 1 0 5256 0 1 4830
box -278 -300 278 300
use sky130_fd_pr__pfet_g5v0d10v5_6ELFTH  XM17
timestamp 1699295625
transform 1 0 4962 0 1 6373
box -308 -339 308 339
use sky130_fd_pr__pfet_g5v0d10v5_6ELFTH  XM18
timestamp 1699295625
transform 1 0 5578 0 1 6373
box -308 -339 308 339
use sky130_fd_pr__nfet_g5v0d10v5_6XHUDR  XM19
timestamp 1699295625
transform 1 0 5256 0 1 4230
box -278 -300 278 300
use sky130_fd_pr__nfet_g5v0d10v5_6XHUDR  XM20
timestamp 1699295625
transform 1 0 4700 0 1 4230
box -278 -300 278 300
use sky130_fd_pr__nfet_g5v0d10v5_6XHUDR  XM21
timestamp 1699295625
transform 1 0 1920 0 1 4230
box -278 -300 278 300
use sky130_fd_pr__pfet_g5v0d10v5_6ELFTH  XM22
timestamp 1699295625
transform 1 0 2498 0 1 6373
box -308 -339 308 339
use sky130_fd_pr__nfet_g5v0d10v5_6XHUDR  XM23
timestamp 1699295625
transform 1 0 1920 0 1 4828
box -278 -300 278 300
use sky130_fd_pr__pfet_g5v0d10v5_6ELFTH  XM24
timestamp 1699295625
transform 1 0 3114 0 1 6373
box -308 -339 308 339
use sky130_fd_pr__pfet_g5v0d10v5_6ELFTH  XM25
timestamp 1699295625
transform 1 0 3730 0 1 6373
box -308 -339 308 339
use sky130_fd_pr__pfet_g5v0d10v5_6ELFTH  XM26
timestamp 1699295625
transform 1 0 4346 0 1 6373
box -308 -339 308 339
use sky130_fd_pr__nfet_g5v0d10v5_6XHUDR  XM27
timestamp 1699295625
transform 1 0 4144 0 1 4230
box -278 -300 278 300
use sky130_fd_pr__nfet_g5v0d10v5_6XHUDR  XM28
timestamp 1699295625
transform 1 0 3588 0 1 4230
box -278 -300 278 300
use sky130_fd_pr__nfet_g5v0d10v5_6XHUDR  XM29
timestamp 1699295625
transform 1 0 3032 0 1 4230
box -278 -300 278 300
use sky130_fd_pr__nfet_g5v0d10v5_6XHUDR  XM30
timestamp 1699295625
transform 1 0 2476 0 1 4230
box -278 -300 278 300
use sky130_fd_pr__pfet_g5v0d10v5_6ELFTH  XM31
timestamp 1699295625
transform 1 0 6194 0 1 5695
box -308 -339 308 339
use sky130_fd_pr__nfet_g5v0d10v5_6XHUDR  XM32
timestamp 1699295625
transform 1 0 5812 0 1 4830
box -278 -300 278 300
use sky130_fd_pr__nfet_g5v0d10v5_6XHUDR  XM33
timestamp 1699295625
transform 1 0 1364 0 1 4828
box -278 -300 278 300
use sky130_fd_pr__pfet_g5v0d10v5_6ELFTH  XM34
timestamp 1699295625
transform 1 0 2498 0 1 5695
box -308 -339 308 339
use sky130_fd_pr__nfet_01v8_L7BSKG  XM35
timestamp 1699295625
transform 1 0 10367 0 1 6113
box -211 -221 211 221
use sky130_fd_pr__nfet_g5v0d10v5_6XHUDR  XM36
timestamp 1699295625
transform 1 0 2476 0 1 4830
box -278 -300 278 300
use sky130_fd_pr__pfet_g5v0d10v5_6ELFTH  XM37
timestamp 1699295625
transform 1 0 6810 0 1 5695
box -308 -339 308 339
use sky130_fd_pr__nfet_g5v0d10v5_6XHUDR  XM38
timestamp 1699295625
transform 1 0 6368 0 1 4830
box -278 -300 278 300
use sky130_fd_pr__pfet_g5v0d10v5_6ELFTH  XM39
timestamp 1699295625
transform 1 0 6194 0 1 6373
box -308 -339 308 339
use sky130_fd_pr__pfet_g5v0d10v5_6ELFTH  XM40
timestamp 1699295625
transform 1 0 6810 0 1 6373
box -308 -339 308 339
use sky130_fd_pr__nfet_g5v0d10v5_6XHUDR  XM41
timestamp 1699295625
transform 1 0 6368 0 1 4230
box -278 -300 278 300
use sky130_fd_pr__nfet_g5v0d10v5_6XHUDR  XM42
timestamp 1699295625
transform 1 0 5812 0 1 4230
box -278 -300 278 300
<< labels >>
flabel metal2 0 7701 200 9695 0 FreeSans 256 0 0 0 avdd
port 0 nsew
flabel metal2 0 1068 200 3062 0 FreeSans 256 0 0 0 avss
port 1 nsew
flabel metal1 12042 3634 12242 4391 0 FreeSans 256 0 0 0 dvdd
port 3 nsew
flabel metal2 12042 4786 12242 4986 0 FreeSans 256 0 0 0 ena
port 4 nsew
flabel metal1 12042 6364 12242 7121 0 FreeSans 256 0 0 0 dvss
port 2 nsew
flabel metal2 12042 5630 12242 5830 0 FreeSans 256 0 0 0 dout
port 5 nsew
flabel metal2 s 12142 7701 12242 9695 0 FreeSans 640 90 0 0 avdd
port 0 nsew
flabel metal2 s 11934 1068 12242 3062 0 FreeSans 960 90 0 0 avss
port 1 nsew
<< properties >>
string FIXED_BBOX 0 0 12242 10724
<< end >>
