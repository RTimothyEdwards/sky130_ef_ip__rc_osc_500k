VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_ef_ip__rc_osc_500k
  CLASS BLOCK ;
  FOREIGN sky130_ef_ip__rc_osc_500k ;
  ORIGIN 0.000 0.000 ;
  SIZE 61.210 BY 53.620 ;
  PIN avdd
    ANTENNADIFFAREA 148.310989 ;
    PORT
      LAYER met2 ;
        RECT 0.000 38.505 60.270 48.475 ;
    END
    PORT
      LAYER met2 ;
        RECT 60.710 38.505 61.210 48.475 ;
    END
  END avdd
  PIN avss
    ANTENNADIFFAREA 114.014595 ;
    PORT
      LAYER met2 ;
        RECT 0.000 5.340 1.595 15.310 ;
    END
    PORT
      LAYER met2 ;
        RECT 59.670 5.340 61.210 15.310 ;
    END
  END avss
  PIN dvss
    ANTENNADIFFAREA 6.628900 ;
    PORT
      LAYER met1 ;
        RECT 59.320 31.820 61.210 35.605 ;
    END
  END dvss
  PIN dvdd
    ANTENNADIFFAREA 4.280700 ;
    PORT
      LAYER met1 ;
        RECT 59.320 18.170 61.210 21.955 ;
    END
  END dvdd
  PIN ena
    ANTENNAGATEAREA 0.858000 ;
    ANTENNADIFFAREA 0.202500 ;
    PORT
      LAYER met2 ;
        RECT 60.210 23.930 61.210 24.930 ;
    END
  END ena
  PIN dout
    ANTENNADIFFAREA 0.556800 ;
    PORT
      LAYER met2 ;
        RECT 60.210 28.150 61.210 29.150 ;
    END
  END dout
  OBS
      LAYER nwell ;
        RECT 0.000 52.010 61.210 53.620 ;
        RECT 0.000 1.610 1.610 52.010 ;
        RECT 0.000 0.000 61.210 1.610 ;
      LAYER li1 ;
        RECT 0.430 0.465 60.755 53.180 ;
      LAYER met1 ;
        RECT 0.430 35.885 60.760 51.000 ;
        RECT 0.430 31.540 59.040 35.885 ;
        RECT 0.430 22.235 60.760 31.540 ;
        RECT 0.430 17.890 59.040 22.235 ;
        RECT 0.430 2.590 60.760 17.890 ;
      LAYER met2 ;
        RECT 0.460 29.430 60.710 38.225 ;
        RECT 0.460 27.870 59.930 29.430 ;
        RECT 0.460 25.210 60.710 27.870 ;
        RECT 0.460 23.650 59.930 25.210 ;
        RECT 0.460 15.590 60.710 23.650 ;
        RECT 1.875 5.340 59.390 15.590 ;
      LAYER met3 ;
        RECT 11.160 13.680 37.435 27.985 ;
      LAYER met4 ;
        RECT 11.555 17.850 37.335 27.990 ;
  END
END sky130_ef_ip__rc_osc_500k
END LIBRARY

