* NGSPICE file created from sky130_ef_ip__rc_osc_500k.ext - technology: sky130A

** x2 ena vdd1v8 vdd3v3 GND GND dout sky130_ef_ip__rc_osc_500k
** .subckt sky130_ef_ip__rc_osc_500k dout dvss dvdd avss avdd ena

.subckt sky130_ef_ip__rc_osc_500k ena dvdd avdd dvss avss dout
X0 a_1178_9768# a_1344_7168# avss.t94 sky130_fd_pr__res_xhigh_po_0p35 l=11
X1 a_10660_3118# a_10494_518# avss.t0 sky130_fd_pr__res_xhigh_po_0p35 l=11
X2 a_4352_3118# a_4186_518# avss.t144 sky130_fd_pr__res_xhigh_po_0p35 l=11
X3 a_6490_9768# a_6656_7168# avss.t138 sky130_fd_pr__res_xhigh_po_0p35 l=11
X4 a_3502_9768# a_3336_7168# avss.t142 sky130_fd_pr__res_xhigh_po_0p35 l=11
X5 a_5162_9768# a_4996_7168# avss.t147 sky130_fd_pr__res_xhigh_po_0p35 l=11
X6 a_8814_9768# a_8648_7168# avss.t93 sky130_fd_pr__res_xhigh_po_0p35 l=11
X7 avdd.t42 a_2858_518# avss.t145 sky130_fd_pr__res_xhigh_po_0p35 l=11
X8 a_7718_4786# ena.t0 a_7560_4786# avss.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X9 a_7154_9768# a_7320_7168# avss.t143 sky130_fd_pr__res_xhigh_po_0p35 l=11
X10 a_5348_3118# a_5182_518# avss.t146 sky130_fd_pr__res_xhigh_po_0p35 l=11
X11 a_11636_7168# a_11490_518# avss.t166 sky130_fd_pr__res_xhigh_po_0p35 l=11
X12 a_4166_9768# a_4000_7168# avss.t56 sky130_fd_pr__res_xhigh_po_0p35 l=11
X13 a_11138_9768# a_11304_7168# avss.t116 sky130_fd_pr__res_xhigh_po_0p35 l=11
X14 a_4194_4788.t0 a_3638_4788.t2 a_4036_4788# avss.t1 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X15 avdd.t31 a_3854_518# avss.t96 sky130_fd_pr__res_xhigh_po_0p35 l=11
X16 a_2506_9768# a_2340_7168# avss.t115 sky130_fd_pr__res_xhigh_po_0p35 l=11
X17 a_9478_9768# a_9312_7168# avss.t68 sky130_fd_pr__res_xhigh_po_0p35 l=11
X18 a_7818_9768# a_7652_7168# avss.t125 sky130_fd_pr__res_xhigh_po_0p35 l=11
X19 a_6344_3118# a_6178_518# avss.t114 sky130_fd_pr__res_xhigh_po_0p35 l=11
X20 avdd.t9 a_2368_4788.t2 a_2368_4788.t3 avdd.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X21 avdd.t8 a_866_518# avss.t45 sky130_fd_pr__res_xhigh_po_0p35 l=11
X22 a_846_9768# a_1012_7168# avss.t55 sky130_fd_pr__res_xhigh_po_0p35 l=11
X23 a_6158_9768# a_6324_7168# avss.t113 sky130_fd_pr__res_xhigh_po_0p35 l=11
X24 a_4684_3118# a_4850_518# avss.t67 sky130_fd_pr__res_xhigh_po_0p35 l=11
X25 a_10806_9768# a_10972_7168# avss.t124 sky130_fd_pr__res_xhigh_po_0p35 l=11
X26 avss.t121 ena.t1 rc_osc_level_shifter_0.outb_h.t1 avss.t120 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X27 a_10142_9768# a_10308_7168# avss.t48 sky130_fd_pr__res_xhigh_po_0p35 l=11
X28 a_7340_3118# a_7174_518# avss.t16 sky130_fd_pr__res_xhigh_po_0p35 l=11
X29 avdd.t30 a_2368_4788.t4 a_4854_5653# avdd.t5 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X30 a_5826_9768# a_5992_7168# avss.t60 sky130_fd_pr__res_xhigh_po_0p35 l=11
X31 a_5162_9768# a_5328_7168# avss.t54 sky130_fd_pr__res_xhigh_po_0p35 l=11
X32 avdd.t45 a_2368_4788.t5 a_5470_5653# avdd.t38 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X33 avdd.t21 a_1862_518# avss.t91 sky130_fd_pr__res_xhigh_po_0p35 l=11
X34 a_5680_3118# a_5846_518# avss.t112 sky130_fd_pr__res_xhigh_po_0p35 l=11
X35 a_9146_9768# a_8980_7168# avss.t15 sky130_fd_pr__res_xhigh_po_0p35 l=11
X36 a_8336_3118# a_8170_518# avss.t90 sky130_fd_pr__res_xhigh_po_0p35 l=11
X37 a_4830_9768# a_4996_7168# avss.t53 sky130_fd_pr__res_xhigh_po_0p35 l=11
X38 avdd.t11 a_2858_518# avss.t52 sky130_fd_pr__res_xhigh_po_0p35 l=11
X39 a_6676_3118# a_6842_518# avss.t111 sky130_fd_pr__res_xhigh_po_0p35 l=11
X40 avdd.t29 a_1530_518# avss.t92 sky130_fd_pr__res_xhigh_po_0p35 l=11
X41 a_10474_9768# a_10640_7168# avss.t51 sky130_fd_pr__res_xhigh_po_0p35 l=11
X42 a_3082_4788.t2 avss.t61 sky130_fd_pr__cap_mim_m3_1 l=6 w=3
X43 a_1842_9768# a_1676_7168# avss.t110 sky130_fd_pr__res_xhigh_po_0p35 l=11
X44 a_9332_3118# a_9166_518# avss.t141 sky130_fd_pr__res_xhigh_po_0p35 l=11
X45 avdd.t39 a_3854_518# avss.t126 sky130_fd_pr__res_xhigh_po_0p35 l=11
X46 avdd.t1 rc_osc_level_shifter_0.out_h.t2 a_2368_4788.t0 avdd.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X47 dvdd.t4 ena.t2 rc_osc_level_shifter_0.inb_l dvdd.t3 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X48 a_5494_9768# a_5660_7168# avss.t36 sky130_fd_pr__res_xhigh_po_0p35 l=11
X49 a_4750_4788.t2 avss.t117 sky130_fd_pr__cap_mim_m3_1 l=6 w=3
X50 a_4750_4788.t1 a_4194_4788.t2 a_4854_5653# avdd.t5 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X51 a_3638_4788.t3 avss.t57 sky130_fd_pr__cap_mim_m3_1 l=6 w=3
X52 a_10328_3118# a_10162_518# avss.t85 sky130_fd_pr__res_xhigh_po_0p35 l=11
X53 a_7672_3118# a_7838_518# avss.t14 sky130_fd_pr__res_xhigh_po_0p35 l=11
X54 a_1414_4786.t3 rc_osc_level_shifter_0.outb_h.t2 avss.t101 avss.t100 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X55 avdd.t40 a_534_518# avss.t130 sky130_fd_pr__res_xhigh_po_0p35 l=11
X56 avdd.t13 a_2526_518# avss.t59 sky130_fd_pr__res_xhigh_po_0p35 l=11
X57 a_1414_4786.t0 rc_osc_level_shifter_0.out_h.t3 a_514_7168.t0 avss.t5 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X58 avdd.t7 a_1198_518# avss.t44 sky130_fd_pr__res_xhigh_po_0p35 l=11
X59 a_5306_4788.t1 a_4750_4788.t3 a_5470_5653# avdd.t38 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X60 a_11324_3118# a_11158_518# avss.t119 sky130_fd_pr__res_xhigh_po_0p35 l=11
X61 a_5016_3118# a_4850_518# avss.t40 sky130_fd_pr__res_xhigh_po_0p35 l=11
X62 a_4498_9768# a_4664_7168# avss.t49 sky130_fd_pr__res_xhigh_po_0p35 l=11
X63 a_5306_4788.t2 avss.t139 sky130_fd_pr__cap_mim_m3_1 l=6 w=3
X64 a_8668_3118# a_8834_518# avss.t136 sky130_fd_pr__res_xhigh_po_0p35 l=11
X65 a_9810_9768# a_9976_7168# avss.t13 sky130_fd_pr__res_xhigh_po_0p35 l=11
X66 avdd.t16 a_2368_4788.t6 a_3622_5653# avdd.t15 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X67 avdd.t35 a_3522_518# avss.t109 sky130_fd_pr__res_xhigh_po_0p35 l=11
X68 avdd.t10 a_2194_518# avss.t50 sky130_fd_pr__res_xhigh_po_0p35 l=11
X69 a_6260_4788# a_1414_4786.t4 avss.t77 avss.t76 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X70 a_3170_9768# a_3004_7168# avss.t135 sky130_fd_pr__res_xhigh_po_0p35 l=11
X71 a_6012_3118# a_5846_518# avss.t89 sky130_fd_pr__res_xhigh_po_0p35 l=11
X72 a_1510_9768# a_1344_7168# avss.t164 sky130_fd_pr__res_xhigh_po_0p35 l=11
X73 a_6822_9768# a_6656_7168# avss.t35 sky130_fd_pr__res_xhigh_po_0p35 l=11
X74 a_8482_9768# a_8316_7168# avss.t129 sky130_fd_pr__res_xhigh_po_0p35 l=11
X75 avdd.t20 a_2368_4788.t7 a_3006_5653# avdd.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X76 a_9664_3118# a_9830_518# avss.t95 sky130_fd_pr__res_xhigh_po_0p35 l=11
X77 avdd.t22 a_2368_4788.t8 a_4238_5653# avdd.t12 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X78 dvss.t5 ena.t3 rc_osc_level_shifter_0.inb_l dvss.t4 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X79 a_10806_9768# a_10640_7168# avss.t165 sky130_fd_pr__res_xhigh_po_0p35 l=11
X80 a_9482_5327# rc_osc_level_shifter_0.out_h.t4 rc_osc_level_shifter_0.outb_h.t0 avdd.t17 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X81 avdd.t33 a_3190_518# avss.t104 sky130_fd_pr__res_xhigh_po_0p35 l=11
X82 a_3502_9768# a_3668_7168# avss.t140 sky130_fd_pr__res_xhigh_po_0p35 l=11
X83 avdd.t24 a_2368_4788.t9 a_6702_5653# avdd.t23 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X84 a_4352_3118# a_4518_518# avss.t39 sky130_fd_pr__res_xhigh_po_0p35 l=11
X85 a_2174_9768# a_2008_7168# avss.t84 sky130_fd_pr__res_xhigh_po_0p35 l=11
X86 a_7486_9768# a_7320_7168# avss.t34 sky130_fd_pr__res_xhigh_po_0p35 l=11
X87 a_10660_3118# a_10826_518# avss.t66 sky130_fd_pr__res_xhigh_po_0p35 l=11
X88 a_5826_9768# a_5660_7168# avss.t83 sky130_fd_pr__res_xhigh_po_0p35 l=11
X89 dout.t2 a_7718_4786# dvdd.t6 dvdd.t5 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X90 a_7008_3118# a_6842_518# avss.t58 sky130_fd_pr__res_xhigh_po_0p35 l=11
X91 avdd.t34 a_1530_518# avss.t108 sky130_fd_pr__res_xhigh_po_0p35 l=11
X92 avdd.t43 a_2368_4788.t10 a_6086_5653# avdd.t37 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X93 a_9332_3118# a_9498_518# avss.t20 sky130_fd_pr__res_xhigh_po_0p35 l=11
X94 a_11890_5939# a_7718_4786# dvss.t7 dvss.t6 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.15
X95 dvss.t3 ena.t4 sky130_fd_pr__diode_pw2nd_05v5 perim=1.8e+06 area=2.025e+11
X96 a_4166_9768# a_4332_7168# avss.t99 sky130_fd_pr__res_xhigh_po_0p35 l=11
X97 a_5348_3118# a_5514_518# avss.t33 sky130_fd_pr__res_xhigh_po_0p35 l=11
X98 avdd.t18 a_4186_518# avss.t79 sky130_fd_pr__res_xhigh_po_0p35 l=11
X99 a_9478_9768# a_9644_7168# avss.t65 sky130_fd_pr__res_xhigh_po_0p35 l=11
X100 a_10328_3118# a_10494_518# avss.t134 sky130_fd_pr__res_xhigh_po_0p35 l=11
X101 a_514_9768# a_680_7168# avss.t38 sky130_fd_pr__res_xhigh_po_0p35 l=11
X102 rc_osc_level_shifter_0.out_h.t1 rc_osc_level_shifter_0.outb_h.t3 a_8714_4659# avdd.t27 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X103 a_1178_9768# a_1012_7168# avss.t32 sky130_fd_pr__res_xhigh_po_0p35 l=11
X104 a_8004_3118# a_7838_518# avss.t133 sky130_fd_pr__res_xhigh_po_0p35 l=11
X105 avdd.t44 a_2526_518# avss.t156 sky130_fd_pr__res_xhigh_po_0p35 l=11
X106 a_5148_4788# a_1414_4786.t5 avss.t75 avss.t74 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X107 a_2982_4700.t0 a_5862_4788# a_6260_4788# avss.t76 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X108 a_8150_9768# a_7984_7168# avss.t64 sky130_fd_pr__res_xhigh_po_0p35 l=11
X109 rc_osc_level_shifter_0.out_h.t0 rc_osc_level_shifter_0.inb_l avss.t42 avss.t41 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X110 a_5704_4788# a_1414_4786.t6 avss.t73 avss.t72 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X111 a_6344_3118# a_6510_518# avss.t132 sky130_fd_pr__res_xhigh_po_0p35 l=11
X112 a_3638_4788.t1 a_3082_4788.t3 a_3622_5653# avdd.t15 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X113 a_11324_3118# a_11490_518# avss.t37 sky130_fd_pr__res_xhigh_po_0p35 l=11
X114 a_5016_3118# a_5182_518# avss.t31 sky130_fd_pr__res_xhigh_po_0p35 l=11
X115 avdd.t19 a_866_518# avss.t88 sky130_fd_pr__res_xhigh_po_0p35 l=11
X116 a_9000_3118# a_8834_518# avss.t155 sky130_fd_pr__res_xhigh_po_0p35 l=11
X117 dvss.t1 rc_osc_level_shifter_0.inb_l dout.t0 dvss.t0 sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.15
X118 a_3480_4788# a_1414_4786.t7 avss.t70 avss.t17 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X119 a_3170_9768# a_3336_7168# avss.t128 sky130_fd_pr__res_xhigh_po_0p35 l=11
X120 a_8482_9768# a_8648_7168# avss.t82 sky130_fd_pr__res_xhigh_po_0p35 l=11
X121 a_3082_4788.t1 a_2982_4700.t2 a_3006_5653# avdd.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X122 a_4194_4788.t1 a_3638_4788.t4 a_4238_5653# avdd.t12 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X123 dvdd.t2 ena.t5 a_7718_4786# dvdd.t1 sky130_fd_pr__pfet_01v8 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.15
X124 a_7154_9768# a_6988_7168# avss.t127 sky130_fd_pr__res_xhigh_po_0p35 l=11
X125 avdd.t6 a_3522_518# avss.t30 sky130_fd_pr__res_xhigh_po_0p35 l=11
X126 a_11138_9768# a_10972_7168# avss.t29 sky130_fd_pr__res_xhigh_po_0p35 l=11
X127 a_2982_4700.t1 a_5862_4788# a_6702_5653# avdd.t23 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X128 a_7340_3118# a_7506_518# avss.t81 sky130_fd_pr__res_xhigh_po_0p35 l=11
X129 a_6012_3118# a_6178_518# avss.t28 sky130_fd_pr__res_xhigh_po_0p35 l=11
X130 a_3834_9768# a_4000_7168# avss.t150 sky130_fd_pr__res_xhigh_po_0p35 l=11
X131 a_9146_9768# a_9312_7168# avss.t87 sky130_fd_pr__res_xhigh_po_0p35 l=11
X132 a_9996_3118# a_9830_518# avss.t154 sky130_fd_pr__res_xhigh_po_0p35 l=11
X133 a_4684_3118# a_4518_518# avss.t163 sky130_fd_pr__res_xhigh_po_0p35 l=11
X134 a_5862_4788# a_5306_4788.t3 a_6086_5653# avdd.t37 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X135 a_10992_3118# a_10826_518# avss.t78 sky130_fd_pr__res_xhigh_po_0p35 l=11
X136 a_8336_3118# a_8502_518# avss.t162 sky130_fd_pr__res_xhigh_po_0p35 l=11
X137 a_6158_9768# a_5992_7168# avss.t153 sky130_fd_pr__res_xhigh_po_0p35 l=11
X138 a_5306_4788.t0 a_4750_4788.t4 a_5148_4788# avss.t74 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X139 a_7008_3118# a_7174_518# avss.t161 sky130_fd_pr__res_xhigh_po_0p35 l=11
X140 a_7718_4786# a_2982_4700.t3 dvdd.t0 avdd.t32 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X141 a_4592_4788# a_1414_4786.t8 avss.t152 avss.t80 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X142 a_5862_4788# a_5306_4788.t4 a_5704_4788# avss.t72 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X143 a_846_9768# a_680_7168# avss.t160 sky130_fd_pr__res_xhigh_po_0p35 l=11
X144 a_8814_9768# a_8980_7168# avss.t159 sky130_fd_pr__res_xhigh_po_0p35 l=11
X145 a_5680_3118# a_5514_518# avss.t71 sky130_fd_pr__res_xhigh_po_0p35 l=11
X146 a_2838_9768# a_3004_7168# avss.t69 sky130_fd_pr__res_xhigh_po_0p35 l=11
X147 avdd.t28 rc_osc_level_shifter_0.out_h.t5 a_8714_4659# avdd.t27 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X148 a_8150_9768# a_8316_7168# avss.t149 sky130_fd_pr__res_xhigh_po_0p35 l=11
X149 a_3638_4788.t0 a_3082_4788.t4 a_3480_4788# avss.t17 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X150 a_2526_4188# a_1414_4786.t9 avss.t22 avss.t21 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X151 a_8004_3118# a_8170_518# avss.t86 sky130_fd_pr__res_xhigh_po_0p35 l=11
X152 a_2924_4788# a_1414_4786.t10 avss.t97 avss.t25 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X153 a_11470_9768# a_11304_7168# avss.t157 sky130_fd_pr__res_xhigh_po_0p35 l=11
X154 a_9482_5327# rc_osc_level_shifter_0.outb_h.t4 avdd.t26 avdd.t25 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X155 a_2506_9768# a_2672_7168# avss.t137 sky130_fd_pr__res_xhigh_po_0p35 l=11
X156 a_7818_9768# a_7984_7168# avss.t19 sky130_fd_pr__res_xhigh_po_0p35 l=11
X157 a_11890_5939# ena.t6 dout.t1 dvss.t2 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.15
X158 a_1842_9768# a_2008_7168# avss.t98 sky130_fd_pr__res_xhigh_po_0p35 l=11
X159 a_6676_3118# a_6510_518# avss.t148 sky130_fd_pr__res_xhigh_po_0p35 l=11
X160 a_6490_9768# a_6324_7168# avss.t12 sky130_fd_pr__res_xhigh_po_0p35 l=11
X161 avdd.t14 a_1198_518# avss.t63 sky130_fd_pr__res_xhigh_po_0p35 l=11
X162 a_4830_9768# a_4664_7168# avss.t151 sky130_fd_pr__res_xhigh_po_0p35 l=11
X163 a_9000_3118# a_9166_518# avss.t158 sky130_fd_pr__res_xhigh_po_0p35 l=11
X164 a_10474_9768# a_10308_7168# avss.t123 sky130_fd_pr__res_xhigh_po_0p35 l=11
X165 a_9996_3118# a_10162_518# avss.t103 sky130_fd_pr__res_xhigh_po_0p35 l=11
X166 a_1510_9768# a_1676_7168# avss.t11 sky130_fd_pr__res_xhigh_po_0p35 l=11
X167 a_4194_4788.t3 avss.t43 sky130_fd_pr__cap_mim_m3_1 l=6 w=3
X168 a_7672_3118# a_7506_518# avss.t10 sky130_fd_pr__res_xhigh_po_0p35 l=11
X169 a_514_9768# a_514_7168.t1 avss.t122 sky130_fd_pr__res_xhigh_po_0p35 l=11
X170 a_6822_9768# a_6988_7168# avss.t102 sky130_fd_pr__res_xhigh_po_0p35 l=11
X171 a_4750_4788.t0 a_4194_4788.t4 a_4592_4788# avss.t80 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X172 avdd.t2 a_2194_518# avss.t9 sky130_fd_pr__res_xhigh_po_0p35 l=11
X173 a_5494_9768# a_5328_7168# avss.t47 sky130_fd_pr__res_xhigh_po_0p35 l=11
X174 a_2526_4188# rc_osc_level_shifter_0.out_h.t6 a_2368_4788.t1 avss.t21 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X175 a_3834_9768# a_3668_7168# avss.t8 sky130_fd_pr__res_xhigh_po_0p35 l=11
X176 a_3082_4788.t0 a_2982_4700.t4 a_2924_4788# avss.t25 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X177 avdd.t36 a_534_518# avss.t118 sky130_fd_pr__res_xhigh_po_0p35 l=11
X178 a_1414_4786.t2 a_1414_4786.t1 avss.t6 avss.t5 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X179 a_7560_4786# a_2982_4700.t5 avss.t24 avss.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X180 a_2174_9768# a_2340_7168# avss.t7 sky130_fd_pr__res_xhigh_po_0p35 l=11
X181 a_7486_9768# a_7652_7168# avss.t46 sky130_fd_pr__res_xhigh_po_0p35 l=11
X182 a_10992_3118# a_11158_518# avss.t4 sky130_fd_pr__res_xhigh_po_0p35 l=11
X183 a_8668_3118# a_8502_518# avss.t3 sky130_fd_pr__res_xhigh_po_0p35 l=11
X184 avdd.t41 a_3190_518# avss.t131 sky130_fd_pr__res_xhigh_po_0p35 l=11
X185 a_4036_4788# a_1414_4786.t11 avss.t2 avss.t1 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X186 a_11470_9768# a_11636_7168# avss.t107 sky130_fd_pr__res_xhigh_po_0p35 l=11
X187 a_2838_9768# a_2672_7168# avss.t106 sky130_fd_pr__res_xhigh_po_0p35 l=11
X188 a_4498_9768# a_4332_7168# avss.t105 sky130_fd_pr__res_xhigh_po_0p35 l=11
X189 a_9810_9768# a_9644_7168# avss.t62 sky130_fd_pr__res_xhigh_po_0p35 l=11
X190 avdd.t3 a_1862_518# avss.t18 sky130_fd_pr__res_xhigh_po_0p35 l=11
X191 a_9664_3118# a_9498_518# avss.t27 sky130_fd_pr__res_xhigh_po_0p35 l=11
X192 a_10142_9768# a_9976_7168# avss.t26 sky130_fd_pr__res_xhigh_po_0p35 l=11
R0 avss.n269 avss.n3 42418.7
R1 avss.n348 avss.n3 42418.7
R2 avss.n348 avss.n4 42418.7
R3 avss.n269 avss.n4 42418.7
R4 avss.n36 avss.n28 42418.7
R5 avss.n322 avss.n28 42418.7
R6 avss.n322 avss.n29 42418.7
R7 avss.n36 avss.n29 42418.7
R8 avss.n300 avss.n299 4540.48
R9 avss.n324 avss.n323 3194
R10 avss.n301 avss.n39 1379.81
R11 avss.n301 avss.n40 1379.81
R12 avss.n314 avss.n40 1379.81
R13 avss.n314 avss.n39 1379.81
R14 avss.n346 avss.n5 1379.81
R15 avss.n346 avss.n6 1379.81
R16 avss.n326 avss.n6 1379.81
R17 avss.n326 avss.n5 1379.81
R18 avss.n331 avss.n22 1379.81
R19 avss.n332 avss.n22 1379.81
R20 avss.n332 avss.n21 1379.81
R21 avss.n331 avss.n21 1379.81
R22 avss.n215 avss.n214 1379.81
R23 avss.n220 avss.n215 1379.81
R24 avss.n221 avss.n220 1379.81
R25 avss.n221 avss.n214 1379.81
R26 avss.n235 avss.n105 1379.81
R27 avss.n234 avss.n105 1379.81
R28 avss.n234 avss.n104 1379.81
R29 avss.n235 avss.n104 1379.81
R30 avss.n240 avss.n98 1379.81
R31 avss.n241 avss.n98 1379.81
R32 avss.n241 avss.n97 1379.81
R33 avss.n240 avss.n97 1379.81
R34 avss.n189 avss.n182 1379.81
R35 avss.n182 avss.n123 1379.81
R36 avss.n178 avss.n123 1379.81
R37 avss.n189 avss.n178 1379.81
R38 avss.n253 avss.n81 1379.81
R39 avss.n252 avss.n81 1379.81
R40 avss.n252 avss.n80 1379.81
R41 avss.n253 avss.n80 1379.81
R42 avss.n258 avss.n74 1379.81
R43 avss.n259 avss.n74 1379.81
R44 avss.n259 avss.n73 1379.81
R45 avss.n258 avss.n73 1379.81
R46 avss.n162 avss.n140 1379.81
R47 avss.n140 avss.n135 1379.81
R48 avss.n136 avss.n135 1379.81
R49 avss.n162 avss.n136 1379.81
R50 avss.n156 avss.n57 1379.81
R51 avss.n156 avss.n58 1379.81
R52 avss.n288 avss.n58 1379.81
R53 avss.n288 avss.n57 1379.81
R54 avss.n290 avss.n49 1379.81
R55 avss.n290 avss.n50 1379.81
R56 avss.n297 avss.n50 1379.81
R57 avss.n297 avss.n49 1379.81
R58 avss.n202 avss.n18 1379.81
R59 avss.n202 avss.n23 1379.81
R60 avss.n217 avss.n23 1379.81
R61 avss.n217 avss.n18 1379.81
R62 avss.n216 avss.n200 1379.81
R63 avss.n216 avss.n208 1379.81
R64 avss.n223 avss.n208 1379.81
R65 avss.n223 avss.n200 1379.81
R66 avss.n209 avss.n106 1379.81
R67 avss.n209 avss.n107 1379.81
R68 avss.n114 avss.n107 1379.81
R69 avss.n114 avss.n106 1379.81
R70 avss.n117 avss.n95 1379.81
R71 avss.n117 avss.n99 1379.81
R72 avss.n179 avss.n99 1379.81
R73 avss.n179 avss.n95 1379.81
R74 avss.n122 avss.n121 1379.81
R75 avss.n190 avss.n121 1379.81
R76 avss.n190 avss.n120 1379.81
R77 avss.n122 avss.n120 1379.81
R78 avss.n175 avss.n82 1379.81
R79 avss.n175 avss.n83 1379.81
R80 avss.n126 avss.n83 1379.81
R81 avss.n126 avss.n82 1379.81
R82 avss.n129 avss.n71 1379.81
R83 avss.n129 avss.n75 1379.81
R84 avss.n137 avss.n75 1379.81
R85 avss.n137 avss.n71 1379.81
R86 avss.n134 avss.n133 1379.81
R87 avss.n163 avss.n133 1379.81
R88 avss.n163 avss.n132 1379.81
R89 avss.n134 avss.n132 1379.81
R90 avss.n152 avss.n62 1379.81
R91 avss.n152 avss.n144 1379.81
R92 avss.n144 avss.n56 1379.81
R93 avss.n62 avss.n56 1379.81
R94 avss.n292 avss.n54 1379.81
R95 avss.n55 avss.n54 1379.81
R96 avss.n55 avss.n48 1379.81
R97 avss.n292 avss.n48 1379.81
R98 avss.n308 avss.n45 1379.81
R99 avss.n310 avss.n44 1379.81
R100 avss.n310 avss.n45 1379.81
R101 avss.t120 avss.n35 934.398
R102 avss.n300 avss.t41 934.398
R103 avss.n321 avss.n30 812.683
R104 avss.n270 avss.n2 804.212
R105 avss.n349 avss.n2 800.46
R106 avss.n31 avss.n30 789.457
R107 avss.n315 avss.n38 697.509
R108 avss.n321 avss.n320 691.125
R109 avss.n271 avss.n268 665.563
R110 avss.n309 avss.n44 562.854
R111 avss.n316 avss.n35 552.742
R112 avss.n319 avss.n31 460.964
R113 avss.n350 avss.n1 360.981
R114 avss.n320 avss.n319 326.962
R115 avss.n267 avss.n1 307.827
R116 avss.n316 avss.n315 236.889
R117 avss.t41 avss.n38 236.889
R118 avss.n64 avss.t24 235.553
R119 avss.n343 avss.t101 234.381
R120 avss.n283 avss.t77 234.012
R121 avss.n264 avss.t73 234.012
R122 avss.n87 avss.t75 234.012
R123 avss.n249 avss.t152 234.012
R124 avss.n246 avss.t2 234.012
R125 avss.n227 avss.t70 234.012
R126 avss.n231 avss.t97 234.012
R127 avss.n337 avss.t22 234.012
R128 avss.n19 avss.t6 233.994
R129 avss.n46 avss.t121 233.939
R130 avss.n33 avss.t42 233.929
R131 avss.t166 avss.t37 213.194
R132 avss.t37 avss.t119 213.194
R133 avss.t119 avss.t4 213.194
R134 avss.t4 avss.t78 213.194
R135 avss.t78 avss.t66 213.194
R136 avss.t66 avss.t0 213.194
R137 avss.t0 avss.t134 213.194
R138 avss.t134 avss.t85 213.194
R139 avss.t85 avss.t103 213.194
R140 avss.t103 avss.t154 213.194
R141 avss.t154 avss.t95 213.194
R142 avss.t157 avss.t107 212.946
R143 avss.t116 avss.t157 212.946
R144 avss.t29 avss.t116 212.946
R145 avss.t124 avss.t29 212.946
R146 avss.t165 avss.t124 212.946
R147 avss.t51 avss.t165 212.946
R148 avss.t123 avss.t51 212.946
R149 avss.t48 avss.t123 212.946
R150 avss.t26 avss.t48 212.946
R151 avss.t13 avss.t26 212.946
R152 avss.t62 avss.t13 212.946
R153 avss.t65 avss.t62 204.929
R154 avss.t95 avss.t27 204.137
R155 avss.n269 avss.t166 202.793
R156 avss.t107 avss.n36 202.572
R157 avss.t68 avss.t65 197.994
R158 avss.t87 avss.t68 197.994
R159 avss.t15 avss.t87 197.994
R160 avss.t159 avss.t15 197.994
R161 avss.t93 avss.t82 197.994
R162 avss.t82 avss.t129 197.994
R163 avss.t129 avss.t149 197.994
R164 avss.t149 avss.t64 197.994
R165 avss.t64 avss.t19 197.994
R166 avss.t19 avss.t125 197.994
R167 avss.t125 avss.t46 197.994
R168 avss.t46 avss.t34 197.994
R169 avss.t34 avss.t143 197.994
R170 avss.t143 avss.t127 197.994
R171 avss.t127 avss.t102 197.964
R172 avss.t102 avss.t35 197.94
R173 avss.t35 avss.t138 197.94
R174 avss.t138 avss.t12 197.94
R175 avss.t12 avss.t113 197.94
R176 avss.t113 avss.t153 197.94
R177 avss.t60 avss.t83 197.94
R178 avss.t83 avss.t36 197.94
R179 avss.t36 avss.t47 197.94
R180 avss.t47 avss.t54 197.94
R181 avss.t54 avss.t147 197.94
R182 avss.t147 avss.t53 197.94
R183 avss.t53 avss.t151 197.94
R184 avss.t151 avss.t49 197.94
R185 avss.t49 avss.t105 197.94
R186 avss.t105 avss.t99 197.94
R187 avss.t99 avss.t56 197.94
R188 avss.t56 avss.t150 197.94
R189 avss.t150 avss.t8 197.94
R190 avss.t8 avss.t140 197.94
R191 avss.t140 avss.t142 197.94
R192 avss.t142 avss.t128 197.94
R193 avss.t128 avss.t135 197.94
R194 avss.t135 avss.t69 197.94
R195 avss.t69 avss.t106 197.94
R196 avss.t106 avss.t137 197.94
R197 avss.t137 avss.t115 197.94
R198 avss.t115 avss.t7 197.94
R199 avss.t7 avss.t84 197.94
R200 avss.t84 avss.t98 197.94
R201 avss.t98 avss.t110 197.94
R202 avss.t110 avss.t11 197.94
R203 avss.t11 avss.t164 197.94
R204 avss.t164 avss.t94 197.94
R205 avss.t32 avss.t55 197.94
R206 avss.t55 avss.t160 197.94
R207 avss.t160 avss.t38 197.94
R208 avss.t38 avss.t122 197.94
R209 avss.t27 avss.t20 191.405
R210 avss.t20 avss.t141 191.405
R211 avss.t141 avss.t158 191.405
R212 avss.t158 avss.t155 191.405
R213 avss.t155 avss.t136 191.405
R214 avss.t136 avss.t3 191.405
R215 avss.t3 avss.t162 191.405
R216 avss.t122 avss.n322 189.195
R217 avss.n38 avss.t159 163.405
R218 avss.n323 avss.t94 146.667
R219 avss.n293 avss.n292 146.25
R220 avss.n292 avss.t23 146.25
R221 avss.n146 avss.n55 146.25
R222 avss.t23 avss.n55 146.25
R223 avss.n285 avss.n62 146.25
R224 avss.t76 avss.n62 146.25
R225 avss.n149 avss.n144 146.25
R226 avss.n144 avss.t76 146.25
R227 avss.n134 avss.n66 146.25
R228 avss.t72 avss.n134 146.25
R229 avss.n164 avss.n163 146.25
R230 avss.n163 avss.t72 146.25
R231 avss.n260 avss.n71 146.25
R232 avss.t74 avss.n71 146.25
R233 avss.n167 avss.n75 146.25
R234 avss.t74 avss.n75 146.25
R235 avss.n251 avss.n82 146.25
R236 avss.t80 avss.n82 146.25
R237 avss.n170 avss.n83 146.25
R238 avss.t80 avss.n83 146.25
R239 avss.n122 avss.n90 146.25
R240 avss.t1 avss.n122 146.25
R241 avss.n191 avss.n190 146.25
R242 avss.n190 avss.t1 146.25
R243 avss.n242 avss.n95 146.25
R244 avss.t17 avss.n95 146.25
R245 avss.n194 avss.n99 146.25
R246 avss.t17 avss.n99 146.25
R247 avss.n233 avss.n106 146.25
R248 avss.t25 avss.n106 146.25
R249 avss.n197 avss.n107 146.25
R250 avss.t25 avss.n107 146.25
R251 avss.n200 avss.n13 146.25
R252 avss.t21 avss.n200 146.25
R253 avss.n208 avss.n207 146.25
R254 avss.t21 avss.n208 146.25
R255 avss.n333 avss.n18 146.25
R256 avss.t5 avss.n18 146.25
R257 avss.n204 avss.n23 146.25
R258 avss.t5 avss.n23 146.25
R259 avss.n295 avss.n49 146.25
R260 avss.t23 avss.n49 146.25
R261 avss.n293 avss.n50 146.25
R262 avss.t23 avss.n50 146.25
R263 avss.n61 avss.n57 146.25
R264 avss.t76 avss.n57 146.25
R265 avss.n285 avss.n58 146.25
R266 avss.t76 avss.n58 146.25
R267 avss.n162 avss.n161 146.25
R268 avss.t72 avss.n162 146.25
R269 avss.n135 avss.n66 146.25
R270 avss.t72 avss.n135 146.25
R271 avss.n258 avss.n257 146.25
R272 avss.t74 avss.n258 146.25
R273 avss.n260 avss.n259 146.25
R274 avss.n259 avss.t74 146.25
R275 avss.n254 avss.n253 146.25
R276 avss.n253 avss.t80 146.25
R277 avss.n252 avss.n251 146.25
R278 avss.t80 avss.n252 146.25
R279 avss.n189 avss.n188 146.25
R280 avss.t1 avss.n189 146.25
R281 avss.n123 avss.n90 146.25
R282 avss.t1 avss.n123 146.25
R283 avss.n240 avss.n239 146.25
R284 avss.t17 avss.n240 146.25
R285 avss.n242 avss.n241 146.25
R286 avss.n241 avss.t17 146.25
R287 avss.n236 avss.n235 146.25
R288 avss.n235 avss.t25 146.25
R289 avss.n234 avss.n233 146.25
R290 avss.t25 avss.n234 146.25
R291 avss.n214 avss.n213 146.25
R292 avss.t21 avss.n214 146.25
R293 avss.n220 avss.n13 146.25
R294 avss.n220 avss.t21 146.25
R295 avss.n331 avss.n330 146.25
R296 avss.t5 avss.n331 146.25
R297 avss.n333 avss.n332 146.25
R298 avss.n332 avss.t5 146.25
R299 avss.n7 avss.n5 146.25
R300 avss.t100 avss.n5 146.25
R301 avss.n8 avss.n6 146.25
R302 avss.t100 avss.n6 146.25
R303 avss.n304 avss.n39 146.25
R304 avss.t41 avss.n39 146.25
R305 avss.n42 avss.n40 146.25
R306 avss.t41 avss.n40 146.25
R307 avss.n311 avss.n310 146.25
R308 avss.n310 avss.t120 146.25
R309 avss.n308 avss.n307 146.25
R310 avss.t86 avss.t133 145.094
R311 avss.t10 avss.t14 145.094
R312 avss.t16 avss.t161 145.094
R313 avss.t161 avss.t58 145.094
R314 avss.t58 avss.t111 145.094
R315 avss.t111 avss.t148 145.094
R316 avss.t114 avss.t132 145.094
R317 avss.t40 avss.t31 145.094
R318 avss.t67 avss.t163 145.094
R319 avss.t131 avss.t109 145.094
R320 avss.t104 avss.t52 145.094
R321 avss.t108 avss.t18 145.094
R322 avss.t92 avss.t63 145.094
R323 avss.t88 avss.t45 145.094
R324 avss.t130 avss.t88 145.094
R325 avss.t118 avss.t130 145.094
R326 avss.n348 avss.t118 142.078
R327 avss.t133 avss.n298 138.101
R328 avss.t162 avss.t90 136.425
R329 avss.t76 avss.t28 135.48
R330 avss.t80 avss.t39 128.487
R331 avss.n153 avss.t112 125.865
R332 avss.t5 avss.t91 124.99
R333 avss.t25 avss.t145 121.495
R334 avss.n177 avss.t79 118.873
R335 avss.t17 avss.t30 117.999
R336 avss.n145 avss.n48 117.207
R337 avss.n298 avss.n48 117.001
R338 avss.n54 avss.n52 117.001
R339 avss.n291 avss.n54 117.001
R340 avss.n59 avss.n56 117.001
R341 avss.n289 avss.n56 117.001
R342 avss.n152 avss.n151 117.001
R343 avss.n155 avss.n152 117.001
R344 avss.n141 avss.n132 117.001
R345 avss.n153 avss.n132 117.001
R346 avss.n133 avss.n68 117.001
R347 avss.n139 avss.n133 117.001
R348 avss.n137 avss.n70 117.001
R349 avss.n138 avss.n137 117.001
R350 avss.n130 avss.n129 117.001
R351 avss.n129 avss.n128 117.001
R352 avss.n126 avss.n124 117.001
R353 avss.n127 avss.n126 117.001
R354 avss.n175 avss.n174 117.001
R355 avss.n176 avss.n175 117.001
R356 avss.n183 avss.n120 117.001
R357 avss.n177 avss.n120 117.001
R358 avss.n121 avss.n92 117.001
R359 avss.n181 avss.n121 117.001
R360 avss.n179 avss.n94 117.001
R361 avss.n180 avss.n179 117.001
R362 avss.n118 avss.n117 117.001
R363 avss.n117 avss.n116 117.001
R364 avss.n114 avss.n112 117.001
R365 avss.n115 avss.n114 117.001
R366 avss.n209 avss.n110 117.001
R367 avss.n210 avss.n209 117.001
R368 avss.n224 avss.n223 117.001
R369 avss.n223 avss.n222 117.001
R370 avss.n216 avss.n15 117.001
R371 avss.n219 avss.n216 117.001
R372 avss.n217 avss.n17 117.001
R373 avss.n218 avss.n217 117.001
R374 avss.n203 avss.n202 117.001
R375 avss.n202 avss.n27 117.001
R376 avss.n297 avss.n296 117.001
R377 avss.n298 avss.n297 117.001
R378 avss.n290 avss.n53 117.001
R379 avss.n291 avss.n290 117.001
R380 avss.n288 avss.n287 117.001
R381 avss.n289 avss.n288 117.001
R382 avss.n157 avss.n156 117.001
R383 avss.n156 avss.n155 117.001
R384 avss.n143 avss.n136 117.001
R385 avss.n153 avss.n136 117.001
R386 avss.n140 avss.n67 117.001
R387 avss.n140 avss.n139 117.001
R388 avss.n73 avss.n69 117.001
R389 avss.n138 avss.n73 117.001
R390 avss.n77 avss.n74 117.001
R391 avss.n128 avss.n74 117.001
R392 avss.n80 avss.n78 117.001
R393 avss.n127 avss.n80 117.001
R394 avss.n85 avss.n81 117.001
R395 avss.n176 avss.n81 117.001
R396 avss.n185 avss.n178 117.001
R397 avss.n178 avss.n177 117.001
R398 avss.n182 avss.n91 117.001
R399 avss.n182 avss.n181 117.001
R400 avss.n97 avss.n93 117.001
R401 avss.n180 avss.n97 117.001
R402 avss.n101 avss.n98 117.001
R403 avss.n116 avss.n98 117.001
R404 avss.n104 avss.n102 117.001
R405 avss.n115 avss.n104 117.001
R406 avss.n109 avss.n105 117.001
R407 avss.n210 avss.n105 117.001
R408 avss.n221 avss.n111 117.001
R409 avss.n222 avss.n221 117.001
R410 avss.n215 avss.n14 117.001
R411 avss.n219 avss.n215 117.001
R412 avss.n21 avss.n16 117.001
R413 avss.n218 avss.n21 117.001
R414 avss.n25 avss.n22 117.001
R415 avss.n27 avss.n22 117.001
R416 avss.n327 avss.n326 117.001
R417 avss.n326 avss.n325 117.001
R418 avss.n346 avss.n345 117.001
R419 avss.n347 avss.n346 117.001
R420 avss.n302 avss.n301 117.001
R421 avss.n301 avss.n300 117.001
R422 avss.n45 avss.n41 117.001
R423 avss.n45 avss.n35 117.001
R424 avss.n314 avss.n313 117.001
R425 avss.n315 avss.n314 117.001
R426 avss.n44 avss.n43 117.001
R427 avss.t9 avss.n219 115.376
R428 avss.t148 avss.n289 113.627
R429 avss.n128 avss.n127 113.627
R430 avss.n116 avss.n115 113.627
R431 avss.n325 avss.n27 113.627
R432 avss.n222 avss.t59 111.879
R433 avss.t23 avss.t81 111.005
R434 avss.t74 avss.t146 111.005
R435 avss.n181 avss.t126 108.383
R436 avss.n299 avss.t90 104.888
R437 avss.n139 avss.t71 101.391
R438 avss.t153 avss.n37 98.9707
R439 avss.n37 avss.t60 98.9707
R440 avss.n204 avss.n203 98.8418
R441 avss.t100 avss.n324 94.3986
R442 avss.t144 avss.n176 87.4061
R443 avss.t72 avss.t71 84.784
R444 avss.t50 avss.n218 83.9099
R445 avss.n294 avss.n52 82.4476
R446 avss.n287 avss.n59 82.0711
R447 avss.n328 avss.n327 82.0711
R448 avss.n327 avss.n26 82.0711
R449 avss.n151 avss.n63 82.0711
R450 avss.n225 avss.n111 82.0711
R451 avss.n225 avss.n224 82.0711
R452 avss.n335 avss.n14 82.0711
R453 avss.n335 avss.n15 82.0711
R454 avss.n108 avss.n102 82.0711
R455 avss.n112 avss.n108 82.0711
R456 avss.n226 avss.n109 82.0711
R457 avss.n226 avss.n110 82.0711
R458 avss.n243 avss.n93 82.0711
R459 avss.n243 avss.n94 82.0711
R460 avss.n113 avss.n101 82.0711
R461 avss.n118 avss.n113 82.0711
R462 avss.n185 avss.n184 82.0711
R463 avss.n184 avss.n183 82.0711
R464 avss.n244 avss.n91 82.0711
R465 avss.n244 avss.n92 82.0711
R466 avss.n84 avss.n78 82.0711
R467 avss.n124 avss.n84 82.0711
R468 avss.n86 avss.n85 82.0711
R469 avss.n174 avss.n86 82.0711
R470 avss.n261 avss.n69 82.0711
R471 avss.n261 avss.n70 82.0711
R472 avss.n125 avss.n77 82.0711
R473 avss.n130 avss.n125 82.0711
R474 avss.n143 avss.n142 82.0711
R475 avss.n142 avss.n141 82.0711
R476 avss.n262 avss.n67 82.0711
R477 avss.n262 avss.n68 82.0711
R478 avss.n157 avss.n63 82.0711
R479 avss.n329 avss.n25 82.0711
R480 avss.n201 avss.n25 82.0711
R481 avss.n24 avss.n16 82.0711
R482 avss.n334 avss.n16 82.0711
R483 avss.n334 avss.n17 82.0711
R484 avss.n203 avss.n201 82.0711
R485 avss.n148 avss.n59 81.6946
R486 avss.n151 avss.n150 81.6946
R487 avss.n211 avss.n111 81.6946
R488 avss.n224 avss.n199 81.6946
R489 avss.n212 avss.n14 81.6946
R490 avss.n206 avss.n15 81.6946
R491 avss.n237 avss.n102 81.6946
R492 avss.n196 avss.n112 81.6946
R493 avss.n109 avss.n103 81.6946
R494 avss.n198 avss.n110 81.6946
R495 avss.n100 avss.n93 81.6946
R496 avss.n193 avss.n94 81.6946
R497 avss.n238 avss.n101 81.6946
R498 avss.n195 avss.n118 81.6946
R499 avss.n186 avss.n185 81.6946
R500 avss.n183 avss.n119 81.6946
R501 avss.n187 avss.n91 81.6946
R502 avss.n192 avss.n92 81.6946
R503 avss.n255 avss.n78 81.6946
R504 avss.n169 avss.n124 81.6946
R505 avss.n85 avss.n79 81.6946
R506 avss.n174 avss.n173 81.6946
R507 avss.n76 avss.n69 81.6946
R508 avss.n166 avss.n70 81.6946
R509 avss.n256 avss.n77 81.6946
R510 avss.n168 avss.n130 81.6946
R511 avss.n159 avss.n143 81.6946
R512 avss.n141 avss.n131 81.6946
R513 avss.n160 avss.n67 81.6946
R514 avss.n165 avss.n68 81.6946
R515 avss.n158 avss.n157 81.6946
R516 avss.n205 avss.n17 81.6946
R517 avss.n147 avss.n52 80.9417
R518 avss.t156 avss.n210 80.4137
R519 avss.n309 avss.n308 78.2942
R520 avss.t1 avss.t126 77.7915
R521 avss.t96 avss.n180 76.9175
R522 avss.n317 avss.n316 75.7785
R523 avss.t81 avss.n291 75.1694
R524 avss.n138 avss.t146 75.1694
R525 avss.t21 avss.t59 74.2953
R526 avss.t45 avss.n347 73.4212
R527 avss.n154 avss.t89 72.5472
R528 avss.n347 avss.t44 71.6731
R529 avss.t21 avss.t9 70.7991
R530 avss.n148 avss.n147 70.3602
R531 avss.n291 avss.t16 69.925
R532 avss.t33 avss.n138 69.925
R533 avss.n180 avss.t30 68.1769
R534 avss.t1 avss.t79 67.3028
R535 avss.n210 avss.t145 64.6807
R536 avss.n218 avss.t91 61.1844
R537 avss.t72 avss.t112 60.3104
R538 avss.t120 avss.n309 59.6593
R539 avss.n176 avss.t39 57.6882
R540 avss.n323 avss.t32 51.2742
R541 avss.n155 avss.t28 50.6958
R542 avss.n311 avss.n43 50.3092
R543 avss.n302 avss.n42 50.106
R544 avss.n139 avss.t33 43.7033
R545 avss.n296 avss.n295 43.1857
R546 avss.n345 avss.n7 41.347
R547 avss.n303 avss.n302 40.4775
R548 avss.n299 avss.t86 40.2071
R549 avss.n146 avss.n145 39.9597
R550 avss.n47 avss.n43 39.8117
R551 avss.n181 avss.t96 36.7109
R552 avss.n38 avss.t93 34.5898
R553 avss.t23 avss.t10 34.0887
R554 avss.t74 avss.t31 34.0887
R555 avss.n222 avss.t156 33.2146
R556 avss.n289 avss.t132 31.4665
R557 avss.t63 avss.t100 30.5925
R558 avss.n219 avss.t50 29.7184
R559 avss.n345 avss.n344 27.9126
R560 avss.t17 avss.t109 27.0962
R561 avss.n177 avss.t144 26.2222
R562 avss.n145 avss.n51 25.3701
R563 avss.n296 avss.n51 25.361
R564 avss.n127 avss.t67 24.4741
R565 avss.n312 avss.n311 23.6684
R566 avss.t25 avss.t52 23.6
R567 avss.n312 avss.n42 23.4269
R568 avss.n155 avss.n154 21.8519
R569 avss.n27 avss.t108 20.9779
R570 avss.t5 avss.t18 20.1038
R571 avss.n324 avss.t44 20.1038
R572 avss.t89 avss.n153 19.2297
R573 avss.n293 avss.n51 17.4857
R574 avss.n115 avss.t104 17.4816
R575 avss.n158 avss.n61 17.1477
R576 avss.n161 avss.n159 17.1477
R577 avss.n161 avss.n160 17.1477
R578 avss.n257 avss.n76 17.1477
R579 avss.n257 avss.n256 17.1477
R580 avss.n255 avss.n254 17.1477
R581 avss.n254 avss.n79 17.1477
R582 avss.n188 avss.n186 17.1477
R583 avss.n188 avss.n187 17.1477
R584 avss.n239 avss.n100 17.1477
R585 avss.n239 avss.n238 17.1477
R586 avss.n237 avss.n236 17.1477
R587 avss.n236 avss.n103 17.1477
R588 avss.n213 avss.n211 17.1477
R589 avss.n213 avss.n212 17.1477
R590 avss.n147 avss.n146 17.1477
R591 avss.n149 avss.n148 17.1477
R592 avss.n150 avss.n149 17.1477
R593 avss.n164 avss.n131 17.1477
R594 avss.n165 avss.n164 17.1477
R595 avss.n167 avss.n166 17.1477
R596 avss.n168 avss.n167 17.1477
R597 avss.n170 avss.n169 17.1477
R598 avss.n191 avss.n119 17.1477
R599 avss.n192 avss.n191 17.1477
R600 avss.n194 avss.n193 17.1477
R601 avss.n195 avss.n194 17.1477
R602 avss.n197 avss.n196 17.1477
R603 avss.n198 avss.n197 17.1477
R604 avss.n207 avss.n199 17.1477
R605 avss.n207 avss.n206 17.1477
R606 avss.n205 avss.n204 17.1477
R607 avss.n328 avss.n7 17.0405
R608 avss.n330 avss.n24 17.0405
R609 avss.n330 avss.n329 17.0405
R610 avss.n26 avss.n8 16.8301
R611 avss.n334 avss.n333 16.8301
R612 avss.n225 avss.n13 16.6249
R613 avss.n233 avss.n108 16.6249
R614 avss.n243 avss.n242 16.6249
R615 avss.n184 avss.n90 16.6249
R616 avss.n251 avss.n84 16.6249
R617 avss.n261 avss.n260 16.6249
R618 avss.n142 avss.n66 16.6249
R619 avss.t80 avss.t163 16.6076
R620 avss.n286 avss.n61 15.7791
R621 avss.n313 avss.n312 15.7042
R622 avss.n295 avss.n294 15.6805
R623 avss.n286 avss.n285 15.2981
R624 avss.n294 avss.n293 15.2981
R625 avss.n307 avss.n306 15.1138
R626 avss.n306 avss.n304 14.9595
R627 avss.n172 avss.n170 14.4911
R628 avss.n116 avss.t131 13.9854
R629 avss.n305 avss.n41 13.6894
R630 avss.n270 avss.n269 12.7179
R631 avss.n36 avss.n31 12.7179
R632 avss.n322 avss.n321 12.7179
R633 avss.n349 avss.n348 12.7179
R634 avss.n344 avss.n8 12.7033
R635 avss.n325 avss.t92 10.4892
R636 avss.n159 avss.n158 10.4659
R637 avss.n160 avss.n76 10.4659
R638 avss.n256 avss.n255 10.4659
R639 avss.n186 avss.n79 10.4659
R640 avss.n187 avss.n100 10.4659
R641 avss.n238 avss.n237 10.4659
R642 avss.n211 avss.n103 10.4659
R643 avss.n150 avss.n131 10.4659
R644 avss.n166 avss.n165 10.4659
R645 avss.n169 avss.n168 10.4659
R646 avss.n173 avss.n119 10.4659
R647 avss.n193 avss.n192 10.4659
R648 avss.n196 avss.n195 10.4659
R649 avss.n199 avss.n198 10.4659
R650 avss.n206 avss.n205 10.4659
R651 avss.n212 avss.n24 10.4574
R652 avss.n329 avss.n328 10.4488
R653 avss.n333 avss.n20 10.4301
R654 avss.n201 avss.n26 10.4152
R655 avss.n335 avss.n334 10.3988
R656 avss.n226 avss.n225 10.3825
R657 avss.n113 avss.n108 10.3825
R658 avss.n244 avss.n243 10.3825
R659 avss.n184 avss.n86 10.3825
R660 avss.n125 avss.n84 10.3825
R661 avss.n262 avss.n261 10.3825
R662 avss.n142 avss.n63 10.3825
R663 avss.n336 avss.n13 10.3029
R664 avss.n233 avss.n232 10.3029
R665 avss.n242 avss.n96 10.3029
R666 avss.n245 avss.n90 10.3029
R667 avss.n251 avss.n250 10.3029
R668 avss.n260 avss.n72 10.3029
R669 avss.n263 avss.n66 10.3029
R670 avss.n285 avss.n284 10.3029
R671 avss.n60 avss.n53 9.81158
R672 avss.n171 avss.n89 9.70903
R673 avss.t76 avss.t114 9.61512
R674 avss.n171 avss.n65 9.37433
R675 avss.n298 avss.t14 6.99295
R676 avss.n128 avss.t40 6.99295
R677 avss.n268 avss.n267 6.53477
R678 avss.n201 avss.n20 6.4005
R679 avss.n336 avss.n335 6.32245
R680 avss.n232 avss.n226 6.32245
R681 avss.n113 avss.n96 6.32245
R682 avss.n245 avss.n244 6.32245
R683 avss.n250 avss.n86 6.32245
R684 avss.n125 avss.n72 6.32245
R685 avss.n263 avss.n262 6.32245
R686 avss.n284 avss.n63 6.32245
R687 avss.n341 avss.n11 6.29691
R688 avss.n287 avss.n60 4.94826
R689 avss.n306 avss.n305 3.79309
R690 avss.n320 avss.n29 3.5246
R691 avss.n37 avss.n29 3.5246
R692 avss.n30 avss.n28 3.5246
R693 avss.n37 avss.n28 3.5246
R694 avss.n4 avss.n2 3.5246
R695 avss.n154 avss.n4 3.5246
R696 avss.n267 avss.n3 3.5246
R697 avss.n154 avss.n3 3.5246
R698 avss.n271 avss.n270 3.07647
R699 avss.n350 avss.n349 2.90959
R700 avss.n173 avss.n172 2.6571
R701 avss.n64 avss.n60 2.3284
R702 avss.n344 avss.n343 2.3255
R703 avss.n47 avss.n46 2.3255
R704 avss.n303 avss.n34 2.3255
R705 avss.n278 avss.n277 2.2484
R706 avss.n10 avss 2.08383
R707 avss.n275 avss.n273 2.06801
R708 avss.n278 avss.n276 2.06752
R709 avss.n307 avss.n47 1.38845
R710 avss.n274 avss.n273 1.25938
R711 avss.n337 avss.n336 1.163
R712 avss.n232 avss.n231 1.163
R713 avss.n227 avss.n96 1.163
R714 avss.n246 avss.n245 1.163
R715 avss.n250 avss.n249 1.163
R716 avss.n87 avss.n72 1.163
R717 avss.n264 avss.n263 1.163
R718 avss.n284 avss.n283 1.163
R719 avss.n20 avss.n19 1.163
R720 avss.n343 avss.n342 1.1255
R721 avss.n305 avss.n32 1.03383
R722 avss.n304 avss.n303 0.925801
R723 avss.n282 avss.n64 0.606932
R724 avss.n229 avss.n1 0.577925
R725 avss.n268 avss.n266 0.577925
R726 avss.n19 avss.n9 0.563
R727 avss.n228 avss.n227 0.563
R728 avss.n231 avss.n230 0.563
R729 avss.n338 avss.n337 0.563
R730 avss.n88 avss.n87 0.563
R731 avss.n249 avss.n248 0.563
R732 avss.n247 avss.n246 0.563
R733 avss.n283 avss.n282 0.563
R734 avss.n265 avss.n264 0.563
R735 avss.n351 avss.n350 0.494944
R736 avss.n272 avss.n271 0.494944
R737 avss.n319 avss.n318 0.4655
R738 avss.n340 avss.n339 0.401201
R739 avss.n281 avss.n272 0.356756
R740 avss.n340 avss.n0 0.304064
R741 avss.n287 avss.n286 0.287571
R742 avss.n342 avss.n9 0.243877
R743 avss.n248 avss.n88 0.230632
R744 avss.n248 avss.n247 0.230632
R745 avss.n247 avss.n89 0.204142
R746 avss.n279 avss.n278 0.181204
R747 avss.n294 avss.n53 0.163374
R748 avss.n280 avss.n12 0.163113
R749 avss.n172 avss.n171 0.143769
R750 avss.n341 avss.n340 0.128227
R751 avss.n313 avss.n41 0.119019
R752 avss avss.n351 0.106457
R753 avss.n88 avss.n65 0.104391
R754 avss.n12 avss.n0 0.0954724
R755 avss.n11 avss.n10 0.068442
R756 avss.n281 avss.n280 0.058173
R757 avss.n46 avss.n32 0.048994
R758 avss.n230 avss.n228 0.0444317
R759 avss.n266 avss.n265 0.0418243
R760 avss.n339 avss.n338 0.0386637
R761 avss.n10 avss 0.0334815
R762 avss.n317 avss.n34 0.0319759
R763 avss.t117 avss.n274 0.0307688
R764 avss.n339 avss.n9 0.0307152
R765 avss.n338 avss.n12 0.0278388
R766 avss.n265 avss.n65 0.0245992
R767 avss.t43 avss.n275 0.0217969
R768 avss.t57 avss.n276 0.0217969
R769 avss.n277 avss.t61 0.0217969
R770 avss.n280 avss.n279 0.0211667
R771 avss.n275 avss.t117 0.0183453
R772 avss.n276 avss.t43 0.0183453
R773 avss.n277 avss.t57 0.0183453
R774 avss.n230 avss.n229 0.0170139
R775 avss.n34 avss.n33 0.0164639
R776 avss.n318 avss.n32 0.0161626
R777 avss.n342 avss.n341 0.0108477
R778 avss.n274 avss.t139 0.0103003
R779 avss.n33 avss.n11 0.0068253
R780 avss.n228 avss.n89 0.00555689
R781 avss.n272 avss 0.00344634
R782 avss.n282 avss.n281 0.00302845
R783 avss.n279 avss.n273 0.000669675
R784 avss.n318 avss.n317 0.000650602
R785 avss.n351 avss.n0 0.000606383
R786 avss.n229 avss.n12 0.000579014
R787 avss.n281 avss.n266 0.000579014
R788 avdd.n268 avdd.n267 32453.4
R789 avdd.n267 avdd.n252 32453.4
R790 avdd.n269 avdd.n268 22625.9
R791 avdd.n321 avdd.n252 22623
R792 avdd.n266 avdd.n250 17294.1
R793 avdd.n266 avdd.n262 17294.1
R794 avdd.n270 avdd.n262 12162.6
R795 avdd.n322 avdd.n250 12161
R796 avdd.n321 avdd.n320 8083.85
R797 avdd.n269 avdd.n253 8069.1
R798 avdd.n320 avdd.n319 6124.84
R799 avdd.n322 avdd.n251 4569.24
R800 avdd.n271 avdd.n270 4561.54
R801 avdd.n271 avdd.n254 3771.24
R802 avdd.n254 avdd.n251 3765.08
R803 avdd.n319 avdd.n253 3546.27
R804 avdd.n265 avdd.n264 1252.21
R805 avdd.n263 avdd.n248 1014.54
R806 avdd.n264 avdd.n261 949.297
R807 avdd.n176 avdd.n166 841.241
R808 avdd.n176 avdd.n167 841.241
R809 avdd.n166 avdd.n165 841.241
R810 avdd.n167 avdd.n165 841.241
R811 avdd.n194 avdd.n142 841.241
R812 avdd.n194 avdd.n143 841.241
R813 avdd.n193 avdd.n143 841.241
R814 avdd.n193 avdd.n142 841.241
R815 avdd.n199 avdd.n136 841.241
R816 avdd.n199 avdd.n137 841.241
R817 avdd.n137 avdd.n135 841.241
R818 avdd.n136 avdd.n135 841.241
R819 avdd.n218 avdd.n109 841.241
R820 avdd.n207 avdd.n109 841.241
R821 avdd.n207 avdd.n110 841.241
R822 avdd.n218 avdd.n110 841.241
R823 avdd.n223 avdd.n105 841.241
R824 avdd.n221 avdd.n105 841.241
R825 avdd.n222 avdd.n221 841.241
R826 avdd.n223 avdd.n222 841.241
R827 avdd.n233 avdd.n43 841.241
R828 avdd.n233 avdd.n44 841.241
R829 avdd.n232 avdd.n44 841.241
R830 avdd.n232 avdd.n43 841.241
R831 avdd.n238 avdd.n39 841.241
R832 avdd.n238 avdd.n40 841.241
R833 avdd.n40 avdd.n33 841.241
R834 avdd.n39 avdd.n33 841.241
R835 avdd.n163 avdd.n161 841.241
R836 avdd.n177 avdd.n161 841.241
R837 avdd.n177 avdd.n160 841.241
R838 avdd.n163 avdd.n160 841.241
R839 avdd.n150 avdd.n145 841.241
R840 avdd.n150 avdd.n146 841.241
R841 avdd.n156 avdd.n146 841.241
R842 avdd.n156 avdd.n145 841.241
R843 avdd.n132 avdd.n131 841.241
R844 avdd.n200 avdd.n132 841.241
R845 avdd.n201 avdd.n200 841.241
R846 avdd.n201 avdd.n131 841.241
R847 avdd.n209 avdd.n121 841.241
R848 avdd.n210 avdd.n209 841.241
R849 avdd.n210 avdd.n108 841.241
R850 avdd.n121 avdd.n108 841.241
R851 avdd.n107 avdd.n103 841.241
R852 avdd.n107 avdd.n104 841.241
R853 avdd.n225 avdd.n104 841.241
R854 avdd.n225 avdd.n103 841.241
R855 avdd.n50 avdd.n46 841.241
R856 avdd.n50 avdd.n47 841.241
R857 avdd.n54 avdd.n47 841.241
R858 avdd.n54 avdd.n46 841.241
R859 avdd.n239 avdd.n35 841.241
R860 avdd.n37 avdd.n35 841.241
R861 avdd.n37 avdd.n34 841.241
R862 avdd.n239 avdd.n34 841.241
R863 avdd.n78 avdd.n71 841.241
R864 avdd.n75 avdd.n71 841.241
R865 avdd.n78 avdd.n70 841.241
R866 avdd.n92 avdd.n65 841.241
R867 avdd.n92 avdd.n66 841.241
R868 avdd.n65 avdd.n64 841.241
R869 avdd.n66 avdd.n64 841.241
R870 avdd.n62 avdd.n59 841.241
R871 avdd.n62 avdd.n60 841.241
R872 avdd.n93 avdd.n60 841.241
R873 avdd.n93 avdd.n59 841.241
R874 avdd.n289 avdd.n287 841.241
R875 avdd.n298 avdd.n287 841.241
R876 avdd.n298 avdd.n292 841.241
R877 avdd.n292 avdd.n289 841.241
R878 avdd.n308 avdd.n279 841.241
R879 avdd.n309 avdd.n279 841.241
R880 avdd.n308 avdd.n280 841.241
R881 avdd.n309 avdd.n280 841.241
R882 avdd.n295 avdd.n256 841.241
R883 avdd.n295 avdd.n257 841.241
R884 avdd.n317 avdd.n257 841.241
R885 avdd.n317 avdd.n256 841.241
R886 avdd.n300 avdd.n282 841.241
R887 avdd.n304 avdd.n282 841.241
R888 avdd.n300 avdd.n283 841.241
R889 avdd.n304 avdd.n283 841.241
R890 avdd.n324 avdd.n248 757.859
R891 avdd.n189 avdd.t1 660.576
R892 avdd.n189 avdd.t9 660.562
R893 avdd.n27 avdd.t24 660.562
R894 avdd.n116 avdd.t22 660.562
R895 avdd.n128 avdd.t16 660.562
R896 avdd.n187 avdd.t20 660.562
R897 avdd.n243 avdd.t45 660.562
R898 avdd.n26 avdd.t43 660.562
R899 avdd.n228 avdd.t30 660.562
R900 avdd.n276 avdd.t26 660.391
R901 avdd.n313 avdd.t28 660.38
R902 avdd.n272 avdd.n261 338.13
R903 avdd.n77 avdd.n61 311.062
R904 avdd.n323 avdd.n249 305.512
R905 avdd.n273 avdd.n272 230.186
R906 avdd.n274 avdd.n260 179.423
R907 avdd.n319 avdd.n318 168.218
R908 avdd.t32 avdd.n77 149.226
R909 avdd.t23 avdd.n61 149.226
R910 avdd.t23 avdd.n63 149.226
R911 avdd.t37 avdd.n36 149.226
R912 avdd.t37 avdd.n38 149.226
R913 avdd.t38 avdd.n45 149.226
R914 avdd.t38 avdd.n48 149.226
R915 avdd.n224 avdd.t5 149.226
R916 avdd.n220 avdd.t5 149.226
R917 avdd.n219 avdd.t12 149.226
R918 avdd.n208 avdd.t12 149.226
R919 avdd.t15 avdd.n123 149.226
R920 avdd.t15 avdd.n134 149.226
R921 avdd.t4 avdd.n144 149.226
R922 avdd.t4 avdd.n147 149.226
R923 avdd.t0 avdd.n162 149.226
R924 avdd.t0 avdd.n164 149.226
R925 avdd.n76 avdd.n70 145.906
R926 avdd.n63 avdd.n36 133.113
R927 avdd.n45 avdd.n38 133.113
R928 avdd.n224 avdd.n48 133.113
R929 avdd.n220 avdd.n219 133.113
R930 avdd.n208 avdd.n123 133.113
R931 avdd.n144 avdd.n134 133.113
R932 avdd.n162 avdd.n147 133.113
R933 avdd.t27 avdd.n281 128.886
R934 avdd.t27 avdd.n284 128.886
R935 avdd.t25 avdd.n255 125.255
R936 avdd.n296 avdd.t17 125.255
R937 avdd.n169 avdd.n159 114.112
R938 avdd.n174 avdd.n169 112.749
R939 avdd.n297 avdd.n281 111.338
R940 avdd.n157 avdd.n148 91.9447
R941 avdd.n203 avdd.n202 91.9447
R942 avdd.n119 avdd.n117 91.9447
R943 avdd.n55 avdd.n29 91.9447
R944 avdd.n56 avdd.n32 91.9447
R945 avdd.n84 avdd.n83 91.9447
R946 avdd.n158 avdd.n153 91.9447
R947 avdd.n227 avdd.n226 91.9447
R948 avdd.n229 avdd.n52 90.0623
R949 avdd.n186 avdd.n140 90.0623
R950 avdd.n204 avdd.n127 90.0623
R951 avdd.n217 avdd.n216 90.0623
R952 avdd.n242 avdd.n28 90.0623
R953 avdd.n87 avdd.n86 90.0623
R954 avdd.n82 avdd.n81 90.0623
R955 avdd.n190 avdd.n152 90.0623
R956 avdd.n191 avdd.n151 85.4593
R957 avdd.n185 avdd.n184 85.4593
R958 avdd.n205 avdd.n122 85.4593
R959 avdd.n215 avdd.n214 85.4593
R960 avdd.n230 avdd.n51 85.4593
R961 avdd.n241 avdd.n31 85.4593
R962 avdd.n80 avdd.n68 85.4593
R963 avdd.n88 avdd.n57 85.4593
R964 avdd.n180 avdd.n151 85.0829
R965 avdd.n182 avdd.n157 85.0829
R966 avdd.n184 avdd.n183 85.0829
R967 avdd.n202 avdd.n130 85.0829
R968 avdd.n122 avdd.n120 85.0829
R969 avdd.n212 avdd.n119 85.0829
R970 avdd.n214 avdd.n213 85.0829
R971 avdd.n101 avdd.n51 85.0829
R972 avdd.n99 avdd.n55 85.0829
R973 avdd.n96 avdd.n56 85.0829
R974 avdd.n98 avdd.n31 85.0829
R975 avdd.n73 avdd.n68 85.0829
R976 avdd.n95 avdd.n57 85.0829
R977 avdd.n83 avdd.n58 85.0829
R978 avdd.n179 avdd.n158 85.0829
R979 avdd.n226 avdd.n102 85.0829
R980 avdd.n191 avdd.n149 83.9534
R981 avdd.n185 avdd.n139 83.9534
R982 avdd.n206 avdd.n205 83.9534
R983 avdd.n215 avdd.n106 83.9534
R984 avdd.n230 avdd.n49 83.9534
R985 avdd.n241 avdd.n30 83.9534
R986 avdd.n89 avdd.n88 83.9534
R987 avdd.n111 avdd.n52 82.824
R988 avdd.n149 avdd.n141 82.824
R989 avdd.n196 avdd.n140 82.824
R990 avdd.n197 avdd.n139 82.824
R991 avdd.n138 avdd.n127 82.824
R992 avdd.n206 avdd.n125 82.824
R993 avdd.n217 avdd.n115 82.824
R994 avdd.n114 avdd.n106 82.824
R995 avdd.n49 avdd.n42 82.824
R996 avdd.n235 avdd.n28 82.824
R997 avdd.n86 avdd.n41 82.824
R998 avdd.n236 avdd.n30 82.824
R999 avdd.n90 avdd.n89 82.824
R1000 avdd.n81 avdd.n67 82.824
R1001 avdd.n168 avdd.n152 82.824
R1002 avdd.n69 avdd.n67 64.4732
R1003 avdd.n288 avdd.n286 51.1301
R1004 avdd.n305 avdd.n303 50.4217
R1005 avdd.n265 avdd.n263 49.7553
R1006 avdd.n79 avdd.n78 46.2505
R1007 avdd.n78 avdd.t32 46.2505
R1008 avdd.n240 avdd.n239 46.2505
R1009 avdd.n239 avdd.t37 46.2505
R1010 avdd.n231 avdd.n46 46.2505
R1011 avdd.t38 avdd.n46 46.2505
R1012 avdd.n103 avdd.n53 46.2505
R1013 avdd.t5 avdd.n103 46.2505
R1014 avdd.n126 avdd.n121 46.2505
R1015 avdd.n121 avdd.t12 46.2505
R1016 avdd.n131 avdd.n129 46.2505
R1017 avdd.t15 avdd.n131 46.2505
R1018 avdd.n192 avdd.n145 46.2505
R1019 avdd.t4 avdd.n145 46.2505
R1020 avdd.n171 avdd.n163 46.2505
R1021 avdd.t0 avdd.n163 46.2505
R1022 avdd.n240 avdd.n33 46.2505
R1023 avdd.t37 avdd.n33 46.2505
R1024 avdd.n232 avdd.n231 46.2505
R1025 avdd.t38 avdd.n232 46.2505
R1026 avdd.n222 avdd.n53 46.2505
R1027 avdd.n222 avdd.t5 46.2505
R1028 avdd.n126 avdd.n110 46.2505
R1029 avdd.n110 avdd.t12 46.2505
R1030 avdd.n135 avdd.n129 46.2505
R1031 avdd.t15 avdd.n135 46.2505
R1032 avdd.n193 avdd.n192 46.2505
R1033 avdd.t4 avdd.n193 46.2505
R1034 avdd.n171 avdd.n165 46.2505
R1035 avdd.t0 avdd.n165 46.2505
R1036 avdd.n85 avdd.n64 46.2505
R1037 avdd.t23 avdd.n64 46.2505
R1038 avdd.n85 avdd.n62 46.2505
R1039 avdd.t23 avdd.n62 46.2505
R1040 avdd.n92 avdd.n91 46.2505
R1041 avdd.t23 avdd.n92 46.2505
R1042 avdd.n238 avdd.n237 46.2505
R1043 avdd.t37 avdd.n238 46.2505
R1044 avdd.n234 avdd.n233 46.2505
R1045 avdd.n233 avdd.t38 46.2505
R1046 avdd.n113 avdd.n105 46.2505
R1047 avdd.n105 avdd.t5 46.2505
R1048 avdd.n124 avdd.n109 46.2505
R1049 avdd.n109 avdd.t12 46.2505
R1050 avdd.n199 avdd.n198 46.2505
R1051 avdd.t15 avdd.n199 46.2505
R1052 avdd.n195 avdd.n194 46.2505
R1053 avdd.n194 avdd.t4 46.2505
R1054 avdd.n176 avdd.n175 46.2505
R1055 avdd.t0 avdd.n176 46.2505
R1056 avdd.n75 avdd.n74 46.2505
R1057 avdd.n94 avdd.n93 46.2505
R1058 avdd.n93 avdd.t23 46.2505
R1059 avdd.n97 avdd.n37 46.2505
R1060 avdd.t37 avdd.n37 46.2505
R1061 avdd.n100 avdd.n47 46.2505
R1062 avdd.t38 avdd.n47 46.2505
R1063 avdd.n118 avdd.n104 46.2505
R1064 avdd.t5 avdd.n104 46.2505
R1065 avdd.n211 avdd.n210 46.2505
R1066 avdd.n210 avdd.t12 46.2505
R1067 avdd.n200 avdd.n133 46.2505
R1068 avdd.n200 avdd.t15 46.2505
R1069 avdd.n181 avdd.n146 46.2505
R1070 avdd.t4 avdd.n146 46.2505
R1071 avdd.n178 avdd.n177 46.2505
R1072 avdd.n177 avdd.t0 46.2505
R1073 avdd.n290 avdd.n256 46.2505
R1074 avdd.t25 avdd.n256 46.2505
R1075 avdd.n259 avdd.n257 46.2505
R1076 avdd.t25 avdd.n257 46.2505
R1077 avdd.n310 avdd.n309 46.2505
R1078 avdd.n309 avdd.t27 46.2505
R1079 avdd.n292 avdd.n291 46.2505
R1080 avdd.t17 avdd.n292 46.2505
R1081 avdd.n303 avdd.n282 46.2505
R1082 avdd.t27 avdd.n282 46.2505
R1083 avdd.n287 avdd.n286 46.2505
R1084 avdd.t17 avdd.n287 46.2505
R1085 avdd.n308 avdd.n307 46.2505
R1086 avdd.t27 avdd.n308 46.2505
R1087 avdd.n307 avdd.n283 46.2505
R1088 avdd.t27 avdd.n283 46.2505
R1089 avdd.n74 avdd.n72 44.9285
R1090 avdd.n0 avdd.t18 42.4171
R1091 avdd.n0 avdd.t39 42.3691
R1092 avdd.n1 avdd.t31 42.3691
R1093 avdd.n2 avdd.t6 42.3691
R1094 avdd.n3 avdd.t35 42.3691
R1095 avdd.n4 avdd.t41 42.3691
R1096 avdd.n5 avdd.t33 42.3691
R1097 avdd.n6 avdd.t11 42.3691
R1098 avdd.n7 avdd.t42 42.3691
R1099 avdd.n8 avdd.t44 42.3691
R1100 avdd.n9 avdd.t13 42.3691
R1101 avdd.n10 avdd.t2 42.3691
R1102 avdd.n11 avdd.t10 42.3691
R1103 avdd.n12 avdd.t21 42.3691
R1104 avdd.n13 avdd.t3 42.3691
R1105 avdd.n14 avdd.t34 42.3691
R1106 avdd.n15 avdd.t29 42.3691
R1107 avdd.n16 avdd.t14 42.3691
R1108 avdd.n17 avdd.t7 42.3691
R1109 avdd.n18 avdd.t8 42.3691
R1110 avdd.n19 avdd.t19 42.3691
R1111 avdd.n20 avdd.t40 42.3691
R1112 avdd.n21 avdd.t36 42.3691
R1113 avdd.n178 avdd.n159 39.8981
R1114 avdd.n72 avdd.n69 39.5797
R1115 avdd.n175 avdd.n174 39.2634
R1116 avdd.n72 avdd.n70 37.0005
R1117 avdd.n71 avdd.n68 37.0005
R1118 avdd.n77 avdd.n71 37.0005
R1119 avdd.n56 avdd.n34 37.0005
R1120 avdd.n36 avdd.n34 37.0005
R1121 avdd.n35 avdd.n31 37.0005
R1122 avdd.n38 avdd.n35 37.0005
R1123 avdd.n55 avdd.n54 37.0005
R1124 avdd.n54 avdd.n45 37.0005
R1125 avdd.n51 avdd.n50 37.0005
R1126 avdd.n50 avdd.n48 37.0005
R1127 avdd.n214 avdd.n107 37.0005
R1128 avdd.n220 avdd.n107 37.0005
R1129 avdd.n119 avdd.n108 37.0005
R1130 avdd.n219 avdd.n108 37.0005
R1131 avdd.n209 avdd.n122 37.0005
R1132 avdd.n209 avdd.n208 37.0005
R1133 avdd.n202 avdd.n201 37.0005
R1134 avdd.n201 avdd.n123 37.0005
R1135 avdd.n184 avdd.n132 37.0005
R1136 avdd.n134 avdd.n132 37.0005
R1137 avdd.n157 avdd.n156 37.0005
R1138 avdd.n156 avdd.n144 37.0005
R1139 avdd.n151 avdd.n150 37.0005
R1140 avdd.n150 avdd.n147 37.0005
R1141 avdd.n170 avdd.n161 37.0005
R1142 avdd.n164 avdd.n161 37.0005
R1143 avdd.n86 avdd.n39 37.0005
R1144 avdd.n39 avdd.n36 37.0005
R1145 avdd.n40 avdd.n30 37.0005
R1146 avdd.n40 avdd.n38 37.0005
R1147 avdd.n43 avdd.n28 37.0005
R1148 avdd.n45 avdd.n43 37.0005
R1149 avdd.n49 avdd.n44 37.0005
R1150 avdd.n48 avdd.n44 37.0005
R1151 avdd.n223 avdd.n52 37.0005
R1152 avdd.n224 avdd.n223 37.0005
R1153 avdd.n221 avdd.n106 37.0005
R1154 avdd.n221 avdd.n220 37.0005
R1155 avdd.n218 avdd.n217 37.0005
R1156 avdd.n219 avdd.n218 37.0005
R1157 avdd.n207 avdd.n206 37.0005
R1158 avdd.n208 avdd.n207 37.0005
R1159 avdd.n136 avdd.n127 37.0005
R1160 avdd.n136 avdd.n123 37.0005
R1161 avdd.n139 avdd.n137 37.0005
R1162 avdd.n137 avdd.n134 37.0005
R1163 avdd.n142 avdd.n140 37.0005
R1164 avdd.n144 avdd.n142 37.0005
R1165 avdd.n149 avdd.n143 37.0005
R1166 avdd.n147 avdd.n143 37.0005
R1167 avdd.n173 avdd.n167 37.0005
R1168 avdd.n167 avdd.n164 37.0005
R1169 avdd.n89 avdd.n66 37.0005
R1170 avdd.n66 avdd.n63 37.0005
R1171 avdd.n60 avdd.n57 37.0005
R1172 avdd.n63 avdd.n60 37.0005
R1173 avdd.n83 avdd.n59 37.0005
R1174 avdd.n61 avdd.n59 37.0005
R1175 avdd.n81 avdd.n65 37.0005
R1176 avdd.n65 avdd.n61 37.0005
R1177 avdd.n166 avdd.n152 37.0005
R1178 avdd.n166 avdd.n162 37.0005
R1179 avdd.n160 avdd.n158 37.0005
R1180 avdd.n162 avdd.n160 37.0005
R1181 avdd.n226 avdd.n225 37.0005
R1182 avdd.n225 avdd.n224 37.0005
R1183 avdd.n317 avdd.n316 37.0005
R1184 avdd.n318 avdd.n317 37.0005
R1185 avdd.n289 avdd.n288 37.0005
R1186 avdd.n289 avdd.n255 37.0005
R1187 avdd.n305 avdd.n304 37.0005
R1188 avdd.n304 avdd.n284 37.0005
R1189 avdd.n299 avdd.n298 37.0005
R1190 avdd.n298 avdd.n297 37.0005
R1191 avdd.n301 avdd.n300 37.0005
R1192 avdd.n300 avdd.n281 37.0005
R1193 avdd.n295 avdd.n294 37.0005
R1194 avdd.n296 avdd.n295 37.0005
R1195 avdd.n294 avdd.n279 37.0005
R1196 avdd.n281 avdd.n279 37.0005
R1197 avdd.n280 avdd.n277 37.0005
R1198 avdd.n284 avdd.n280 37.0005
R1199 avdd.n76 avdd.n75 36.2372
R1200 avdd.n73 avdd.n58 35.7439
R1201 avdd.n319 avdd.n254 35.604
R1202 avdd.n311 avdd.n310 26.6196
R1203 avdd.n315 avdd.n259 25.9151
R1204 avdd.n260 avdd.n249 25.2054
R1205 avdd.n82 avdd.n80 24.1639
R1206 avdd.n172 avdd.n170 24.0137
R1207 avdd.n173 avdd.n172 23.5906
R1208 avdd.n303 avdd.n302 23.2301
R1209 avdd.n302 avdd.n286 23.2301
R1210 avdd.n316 avdd.n258 23.1206
R1211 avdd.n316 avdd.n315 23.0608
R1212 avdd.n306 avdd.n305 23.0608
R1213 avdd.n306 avdd.n277 23.0608
R1214 avdd.n288 avdd.n258 22.7005
R1215 avdd.n311 avdd.n277 21.9434
R1216 avdd.n310 avdd.n278 20.2328
R1217 avdd.n278 avdd.n259 20.2328
R1218 avdd.n294 avdd.n285 19.0862
R1219 avdd.n91 avdd.n67 17.1477
R1220 avdd.n91 avdd.n90 17.1477
R1221 avdd.n237 avdd.n41 17.1477
R1222 avdd.n237 avdd.n236 17.1477
R1223 avdd.n235 avdd.n234 17.1477
R1224 avdd.n234 avdd.n42 17.1477
R1225 avdd.n114 avdd.n113 17.1477
R1226 avdd.n124 avdd.n115 17.1477
R1227 avdd.n125 avdd.n124 17.1477
R1228 avdd.n198 avdd.n138 17.1477
R1229 avdd.n198 avdd.n197 17.1477
R1230 avdd.n196 avdd.n195 17.1477
R1231 avdd.n195 avdd.n141 17.1477
R1232 avdd.n175 avdd.n168 17.1477
R1233 avdd.n74 avdd.n73 17.1477
R1234 avdd.n94 avdd.n58 17.1477
R1235 avdd.n95 avdd.n94 17.1477
R1236 avdd.n97 avdd.n96 17.1477
R1237 avdd.n98 avdd.n97 17.1477
R1238 avdd.n100 avdd.n99 17.1477
R1239 avdd.n101 avdd.n100 17.1477
R1240 avdd.n118 avdd.n102 17.1477
R1241 avdd.n213 avdd.n118 17.1477
R1242 avdd.n212 avdd.n211 17.1477
R1243 avdd.n211 avdd.n120 17.1477
R1244 avdd.n133 avdd.n130 17.1477
R1245 avdd.n183 avdd.n133 17.1477
R1246 avdd.n182 avdd.n181 17.1477
R1247 avdd.n181 avdd.n180 17.1477
R1248 avdd.n179 avdd.n178 17.1477
R1249 avdd.n302 avdd.n301 16.2647
R1250 avdd.n90 avdd.n41 15.2961
R1251 avdd.n236 avdd.n235 15.2961
R1252 avdd.n111 avdd.n42 15.2961
R1253 avdd.n115 avdd.n114 15.2961
R1254 avdd.n138 avdd.n125 15.2961
R1255 avdd.n197 avdd.n196 15.2961
R1256 avdd.n168 avdd.n141 15.2961
R1257 avdd.n96 avdd.n95 15.2961
R1258 avdd.n99 avdd.n98 15.2961
R1259 avdd.n102 avdd.n101 15.2961
R1260 avdd.n213 avdd.n212 15.2961
R1261 avdd.n130 avdd.n120 15.2961
R1262 avdd.n183 avdd.n182 15.2961
R1263 avdd.n180 avdd.n179 15.2961
R1264 avdd.n290 avdd.n258 15.193
R1265 avdd.n307 avdd.n306 14.8746
R1266 avdd.n172 avdd.n171 14.4286
R1267 avdd.n299 avdd.n285 13.2702
R1268 avdd.n192 avdd.n191 11.9584
R1269 avdd.n185 avdd.n129 11.9584
R1270 avdd.n205 avdd.n126 11.9584
R1271 avdd.n215 avdd.n53 11.9584
R1272 avdd.n231 avdd.n230 11.9584
R1273 avdd.n241 avdd.n240 11.9584
R1274 avdd.n88 avdd.n85 11.9584
R1275 avdd.n80 avdd.n79 11.9302
R1276 avdd.n307 avdd.n285 11.6153
R1277 avdd.n291 avdd.n285 11.365
R1278 avdd.n112 avdd.n111 10.8684
R1279 avdd.n191 avdd.n190 9.77806
R1280 avdd.n186 avdd.n185 9.77806
R1281 avdd.n205 avdd.n204 9.77806
R1282 avdd.n216 avdd.n215 9.77806
R1283 avdd.n230 avdd.n229 9.77806
R1284 avdd.n242 avdd.n241 9.77806
R1285 avdd.n88 avdd.n87 9.77806
R1286 avdd.n294 avdd.n293 8.8005
R1287 avdd.n170 avdd.n159 8.25174
R1288 avdd.n174 avdd.n173 8.14595
R1289 avdd.t32 avdd.n76 8.02261
R1290 avdd.n293 avdd.n278 7.6005
R1291 avdd.n113 avdd.n112 6.27974
R1292 avdd.n272 avdd.n271 6.16717
R1293 avdd.n271 avdd.n253 6.16717
R1294 avdd.n251 avdd.n249 6.16717
R1295 avdd.n320 avdd.n251 6.16717
R1296 avdd.n273 avdd.n254 4.74409
R1297 avdd.n318 avdd.n255 3.63107
R1298 avdd.t17 avdd.t25 3.63107
R1299 avdd.n297 avdd.n296 3.63107
R1300 avdd.n172 avdd.n169 3.36892
R1301 avdd.n270 avdd.n261 3.36414
R1302 avdd.n270 avdd.n269 3.36414
R1303 avdd.n323 avdd.n322 3.36414
R1304 avdd.n322 avdd.n321 3.36414
R1305 avdd.n312 avdd.n311 3.10844
R1306 avdd.n315 avdd.n314 3.1005
R1307 avdd.n274 avdd.n273 2.57768
R1308 avdd.n79 avdd.n69 2.51578
R1309 avdd.n22 avdd.n21 1.46517
R1310 avdd.n275 avdd.n247 1.34749
R1311 avdd.n266 avdd.n265 1.20965
R1312 avdd.n267 avdd.n266 1.20965
R1313 avdd.n264 avdd.n262 1.05164
R1314 avdd.n268 avdd.n262 1.05164
R1315 avdd.n250 avdd.n248 1.05164
R1316 avdd.n252 avdd.n250 1.05164
R1317 avdd.n293 avdd.n276 0.9305
R1318 avdd.n314 avdd.n275 0.877364
R1319 avdd.n329 avdd.n22 0.87315
R1320 avdd.n187 avdd.n186 0.7755
R1321 avdd.n204 avdd.n128 0.7755
R1322 avdd.n216 avdd.n116 0.7755
R1323 avdd.n243 avdd.n242 0.7755
R1324 avdd.n87 avdd.n26 0.7755
R1325 avdd.n82 avdd.n27 0.7755
R1326 avdd.n190 avdd.n189 0.7755
R1327 avdd.n229 avdd.n228 0.7755
R1328 avdd.n324 avdd.n323 0.621859
R1329 avdd.n24 avdd.n23 0.552286
R1330 avdd.n260 avdd.n247 0.504
R1331 avdd.n325 avdd.n324 0.490106
R1332 avdd.n228 avdd.n25 0.3755
R1333 avdd.n154 avdd.n116 0.3755
R1334 avdd.n188 avdd.n128 0.3755
R1335 avdd.n188 avdd.n187 0.3755
R1336 avdd.n189 avdd.n188 0.3755
R1337 avdd.n244 avdd.n27 0.3755
R1338 avdd.n244 avdd.n26 0.3755
R1339 avdd.n244 avdd.n243 0.3755
R1340 avdd.n291 avdd.n290 0.359379
R1341 avdd.n171 avdd.n153 0.281202
R1342 avdd.n192 avdd.n148 0.281202
R1343 avdd.n203 avdd.n129 0.281202
R1344 avdd.n126 avdd.n117 0.281202
R1345 avdd.n227 avdd.n53 0.281202
R1346 avdd.n231 avdd.n29 0.281202
R1347 avdd.n240 avdd.n32 0.281202
R1348 avdd.n85 avdd.n84 0.281202
R1349 avdd.n327 avdd.n326 0.27802
R1350 avdd.n263 avdd.n22 0.2618
R1351 avdd.n326 avdd.n247 0.244654
R1352 avdd.n154 avdd.n25 0.244171
R1353 avdd.n275 avdd.n274 0.233
R1354 avdd.n246 avdd.n24 0.221333
R1355 avdd.n329 avdd.n328 0.192137
R1356 avdd.n328 avdd.n327 0.185806
R1357 avdd.n112 avdd.n24 0.172219
R1358 avdd.n155 avdd.n154 0.14963
R1359 avdd.n314 avdd.n313 0.122295
R1360 avdd.n245 avdd.n25 0.121149
R1361 avdd.n313 avdd.n312 0.119303
R1362 avdd.n301 avdd.n299 0.117931
R1363 avdd.n326 avdd.n325 0.090332
R1364 avdd.n328 avdd.n23 0.0714439
R1365 avdd.n327 avdd.n246 0.0714439
R1366 avdd.n186 avdd.n148 0.0573889
R1367 avdd.n204 avdd.n203 0.0573889
R1368 avdd.n216 avdd.n117 0.0573889
R1369 avdd.n242 avdd.n29 0.0573889
R1370 avdd.n87 avdd.n32 0.0573889
R1371 avdd.n84 avdd.n82 0.0573889
R1372 avdd.n190 avdd.n153 0.0573889
R1373 avdd.n229 avdd.n227 0.0573889
R1374 avdd.n155 avdd.n23 0.0547069
R1375 avdd.n246 avdd.n245 0.0547069
R1376 avdd.n1 avdd.n0 0.0485324
R1377 avdd.n2 avdd.n1 0.0485324
R1378 avdd.n3 avdd.n2 0.0485324
R1379 avdd.n4 avdd.n3 0.0485324
R1380 avdd.n5 avdd.n4 0.0485324
R1381 avdd.n6 avdd.n5 0.0485324
R1382 avdd.n7 avdd.n6 0.0485324
R1383 avdd.n8 avdd.n7 0.0485324
R1384 avdd.n9 avdd.n8 0.0485324
R1385 avdd.n10 avdd.n9 0.0485324
R1386 avdd.n11 avdd.n10 0.0485324
R1387 avdd.n12 avdd.n11 0.0485324
R1388 avdd.n13 avdd.n12 0.0485324
R1389 avdd.n14 avdd.n13 0.0485324
R1390 avdd.n15 avdd.n14 0.0485324
R1391 avdd.n16 avdd.n15 0.0485324
R1392 avdd.n17 avdd.n16 0.0485324
R1393 avdd.n18 avdd.n17 0.0485324
R1394 avdd.n19 avdd.n18 0.0485324
R1395 avdd.n20 avdd.n19 0.0485324
R1396 avdd.n21 avdd.n20 0.0485324
R1397 avdd avdd.n329 0.0146048
R1398 avdd.n312 avdd 0.0139615
R1399 avdd.n313 avdd.n276 0.00377715
R1400 avdd.n325 avdd 0.00325827
R1401 avdd.n188 avdd.n155 0.000801568
R1402 avdd.n245 avdd.n244 0.000801568
R1403 ena.n5 ena.t2 396.2
R1404 ena.n5 ena.t3 381.825
R1405 ena.n1 ena.t5 305.348
R1406 ena.n0 ena.t6 302.945
R1407 ena.n3 ena.t4 196.596
R1408 ena.n2 ena.t0 112.272
R1409 ena.n2 ena.t1 110.207
R1410 ena.n5 ena.n4 4.5005
R1411 ena.n4 ena.n3 2.03668
R1412 ena.n4 ena.n1 1.72267
R1413 ena.n3 ena.n2 1.20571
R1414 ena.n1 ena.n0 1.06763
R1415 ena.n0 ena 0.368556
R1416 ena ena.n5 0.062375
R1417 a_3638_4788.t1 a_3638_4788.t3 660.754
R1418 a_3638_4788.t3 a_3638_4788.t0 235.388
R1419 a_3638_4788.t3 a_3638_4788.t4 107.769
R1420 a_3638_4788.t3 a_3638_4788.t2 105.281
R1421 a_4194_4788.t1 a_4194_4788.t3 660.745
R1422 a_4194_4788.t3 a_4194_4788.t0 235.613
R1423 a_4194_4788.t3 a_4194_4788.t2 107.96
R1424 a_4194_4788.t3 a_4194_4788.t4 105.281
R1425 a_2368_4788.n1 a_2368_4788.t0 660.24
R1426 a_2368_4788.t3 a_2368_4788.n1 660.24
R1427 a_2368_4788.n1 a_2368_4788.t1 236.429
R1428 a_2368_4788.n0 a_2368_4788.t9 107.941
R1429 a_2368_4788.n1 a_2368_4788.t2 106.373
R1430 a_2368_4788.n0 a_2368_4788.t7 106.373
R1431 a_2368_4788.n0 a_2368_4788.t6 106.373
R1432 a_2368_4788.n0 a_2368_4788.t8 106.373
R1433 a_2368_4788.n0 a_2368_4788.t4 106.373
R1434 a_2368_4788.n0 a_2368_4788.t5 106.373
R1435 a_2368_4788.n0 a_2368_4788.t10 106.373
R1436 a_2368_4788.n1 a_2368_4788.n0 11.6107
R1437 rc_osc_level_shifter_0.outb_h.n0 rc_osc_level_shifter_0.outb_h.t0 660.24
R1438 rc_osc_level_shifter_0.outb_h.n0 rc_osc_level_shifter_0.outb_h.t1 235.004
R1439 rc_osc_level_shifter_0.outb_h rc_osc_level_shifter_0.outb_h.t2 127.82
R1440 rc_osc_level_shifter_0.outb_h.n0 rc_osc_level_shifter_0.outb_h.t3 116.334
R1441 rc_osc_level_shifter_0.outb_h.n0 rc_osc_level_shifter_0.outb_h.t4 107.222
R1442 rc_osc_level_shifter_0.outb_h rc_osc_level_shifter_0.outb_h.n0 11.5134
R1443 a_3082_4788.t1 a_3082_4788.t2 660.769
R1444 a_3082_4788.t2 a_3082_4788.t0 235.127
R1445 a_3082_4788.t2 a_3082_4788.t3 107.582
R1446 a_3082_4788.t2 a_3082_4788.t4 105.273
R1447 rc_osc_level_shifter_0.out_h rc_osc_level_shifter_0.out_h.t1 660.24
R1448 rc_osc_level_shifter_0.out_h rc_osc_level_shifter_0.out_h.t0 235.251
R1449 rc_osc_level_shifter_0.out_h rc_osc_level_shifter_0.out_h.t4 116.338
R1450 rc_osc_level_shifter_0.out_h.n0 rc_osc_level_shifter_0.out_h.t2 110.648
R1451 rc_osc_level_shifter_0.out_h rc_osc_level_shifter_0.out_h.t5 106.773
R1452 rc_osc_level_shifter_0.out_h.n0 rc_osc_level_shifter_0.out_h.t6 106.382
R1453 rc_osc_level_shifter_0.out_h.n0 rc_osc_level_shifter_0.out_h.t3 104.746
R1454 rc_osc_level_shifter_0.out_h rc_osc_level_shifter_0.out_h.n0 21.9372
R1455 dvdd.n18 dvdd.n13 1312.94
R1456 dvdd.n22 dvdd.n12 1312.94
R1457 dvdd.n22 dvdd.n13 1312.94
R1458 dvdd.n5 dvdd.n4 1312.94
R1459 dvdd.n26 dvdd.n25 1108.24
R1460 dvdd.n25 dvdd.n8 1108.24
R1461 dvdd.n6 dvdd.n5 704.168
R1462 dvdd.n34 dvdd.n3 697.11
R1463 dvdd.n37 dvdd.t0 668.082
R1464 dvdd.n0 dvdd.t2 662.312
R1465 dvdd.n31 dvdd.n3 596.572
R1466 dvdd.n31 dvdd.n6 589.715
R1467 dvdd.n26 dvdd.n6 497.647
R1468 dvdd.n8 dvdd.n3 497.647
R1469 dvdd.n24 dvdd.n23 345.777
R1470 dvdd.n32 dvdd.t1 334.182
R1471 dvdd.n24 dvdd.t1 332.08
R1472 dvdd.t3 dvdd.n32 332.08
R1473 dvdd.n33 dvdd.n4 277.072
R1474 dvdd.n23 dvdd.t5 264.262
R1475 dvdd.n18 dvdd.n17 237.584
R1476 dvdd.n39 dvdd.t4 228.498
R1477 dvdd.n9 dvdd.t6 228.239
R1478 dvdd.n20 dvdd.n19 137.024
R1479 dvdd.t3 dvdd.n5 106.007
R1480 dvdd.n19 dvdd.n16 100.001
R1481 dvdd.n20 dvdd.n12 95.2318
R1482 dvdd.n16 dvdd.n13 92.5005
R1483 dvdd.n13 dvdd.t5 92.5005
R1484 dvdd.n27 dvdd.n26 92.5005
R1485 dvdd.n26 dvdd.t1 92.5005
R1486 dvdd.n35 dvdd.n34 92.5005
R1487 dvdd.n28 dvdd.n5 92.5005
R1488 dvdd.n14 dvdd.n8 92.5005
R1489 dvdd.n8 dvdd.t1 92.5005
R1490 dvdd.n28 dvdd.n2 90.9905
R1491 dvdd.n29 dvdd.n28 75.1118
R1492 dvdd.n34 dvdd.n33 74.3381
R1493 dvdd.n17 dvdd.n12 70.7763
R1494 dvdd.n30 dvdd.n29 62.9034
R1495 dvdd.n25 dvdd.n11 61.6672
R1496 dvdd.n25 dvdd.n24 61.6672
R1497 dvdd.n30 dvdd.n1 57.4176
R1498 dvdd.n27 dvdd.n7 53.0829
R1499 dvdd.n29 dvdd.n27 53.0829
R1500 dvdd.n35 dvdd.n2 52.7584
R1501 dvdd.n19 dvdd.n18 46.2505
R1502 dvdd.n4 dvdd.n2 46.2505
R1503 dvdd.n31 dvdd.n30 46.2505
R1504 dvdd.n32 dvdd.n31 46.2505
R1505 dvdd.n22 dvdd.n21 46.2505
R1506 dvdd.n23 dvdd.n22 46.2505
R1507 dvdd.n21 dvdd.n20 44.1706
R1508 dvdd.n15 dvdd.n14 40.0601
R1509 dvdd.n16 dvdd.n15 23.8938
R1510 dvdd.n33 dvdd.t3 21.4216
R1511 dvdd.n17 dvdd.t5 16.7394
R1512 dvdd.n36 dvdd.n1 13.4634
R1513 dvdd.n14 dvdd.n1 12.4864
R1514 dvdd.n11 dvdd.n10 9.51845
R1515 dvdd.n15 dvdd.n11 3.41383
R1516 dvdd.n37 dvdd.n36 2.3255
R1517 dvdd.n10 dvdd.n7 1.83845
R1518 dvdd.n10 dvdd.n9 1.55446
R1519 dvdd.n21 dvdd.n7 0.459987
R1520 dvdd.n39 dvdd.n38 0.317167
R1521 dvdd.n40 dvdd.n39 0.153726
R1522 dvdd.n40 dvdd.n0 0.146137
R1523 dvdd.n36 dvdd.n35 0.129793
R1524 dvdd.n9 dvdd.n0 0.0618011
R1525 dvdd.n38 dvdd.n37 0.038
R1526 dvdd.n41 dvdd.n40 0.0228214
R1527 dvdd dvdd.n41 0.0228214
R1528 dvdd.n38 dvdd 0.004875
R1529 dvdd.n41 dvdd 0.001125
R1530 a_4750_4788.t1 a_4750_4788.t2 660.756
R1531 a_4750_4788.t2 a_4750_4788.t0 235.773
R1532 a_4750_4788.t2 a_4750_4788.t3 108.153
R1533 a_4750_4788.t2 a_4750_4788.t4 105.281
R1534 a_1414_4786.n0 a_1414_4786.t3 237.433
R1535 a_1414_4786.t0 a_1414_4786.n0 235.407
R1536 a_1414_4786.n0 a_1414_4786.t2 233.657
R1537 a_1414_4786.n0 a_1414_4786.t10 113.971
R1538 a_1414_4786.n0 a_1414_4786.t4 105.537
R1539 a_1414_4786.n0 a_1414_4786.t1 104.177
R1540 a_1414_4786.n0 a_1414_4786.t6 104.175
R1541 a_1414_4786.n0 a_1414_4786.t5 104.175
R1542 a_1414_4786.n0 a_1414_4786.t8 104.175
R1543 a_1414_4786.n0 a_1414_4786.t11 104.175
R1544 a_1414_4786.n0 a_1414_4786.t7 104.175
R1545 a_1414_4786.n0 a_1414_4786.t9 104.175
R1546 a_514_7168.t1 a_514_7168.t0 245.28
R1547 a_5306_4788.t1 a_5306_4788.t2 660.806
R1548 a_5306_4788.t2 a_5306_4788.t0 235.982
R1549 a_5306_4788.t2 a_5306_4788.t3 108.346
R1550 a_5306_4788.t2 a_5306_4788.t4 105.281
R1551 dvss.n42 dvss.n38 25476.2
R1552 dvss.n43 dvss.n19 9928.12
R1553 dvss.n62 dvss.n11 2126.44
R1554 dvss.n24 dvss.n11 2126.44
R1555 dvss.n62 dvss.n12 2126.44
R1556 dvss.n24 dvss.n12 2126.44
R1557 dvss.n40 dvss.n35 1836.74
R1558 dvss.n44 dvss.n35 1836.74
R1559 dvss.n44 dvss.n34 1836.74
R1560 dvss.n37 dvss.n9 1836.74
R1561 dvss.n65 dvss.n9 1836.74
R1562 dvss.n37 dvss.n10 1836.74
R1563 dvss.n65 dvss.n10 1836.74
R1564 dvss.n54 dvss.n22 1790.38
R1565 dvss.n22 dvss.n20 1790.38
R1566 dvss.n21 dvss.n20 1790.38
R1567 dvss.n54 dvss.n21 1790.38
R1568 dvss.n64 dvss.n63 1740.52
R1569 dvss.n25 dvss.n23 1449.84
R1570 dvss.n56 dvss.n17 1407.97
R1571 dvss.n56 dvss.n18 1407.97
R1572 dvss.n49 dvss.n17 1407.97
R1573 dvss.n49 dvss.n18 1407.97
R1574 dvss.t2 dvss.n43 818.846
R1575 dvss.n41 dvss.n40 776.158
R1576 dvss.n38 dvss.t6 667.819
R1577 dvss.n64 dvss.t6 667.819
R1578 dvss.n27 dvss.n26 592.715
R1579 dvss.n63 dvss.t4 569.837
R1580 dvss.n48 dvss.t3 468.853
R1581 dvss.n55 dvss.t0 367.87
R1582 dvss.n42 dvss.n41 329.875
R1583 dvss.n26 dvss.t4 317.377
R1584 dvss.n41 dvss.n34 316.318
R1585 dvss.n13 dvss.n11 294.214
R1586 dvss.n10 dvss.n8 292.5
R1587 dvss.t6 dvss.n10 292.5
R1588 dvss.n9 dvss.n7 292.5
R1589 dvss.t6 dvss.n9 292.5
R1590 dvss.n40 dvss.n39 292.5
R1591 dvss.n45 dvss.n44 292.5
R1592 dvss.n44 dvss.t2 292.5
R1593 dvss.n18 dvss.n15 292.5
R1594 dvss.t3 dvss.n18 292.5
R1595 dvss.n54 dvss.n53 292.5
R1596 dvss.t0 dvss.n54 292.5
R1597 dvss.n50 dvss.n49 292.5
R1598 dvss.n49 dvss.n48 292.5
R1599 dvss.n31 dvss.n17 292.5
R1600 dvss.t3 dvss.n17 292.5
R1601 dvss.n30 dvss.n20 292.5
R1602 dvss.t0 dvss.n20 292.5
R1603 dvss.n57 dvss.n56 292.5
R1604 dvss.n56 dvss.n55 292.5
R1605 dvss.n60 dvss.n12 292.5
R1606 dvss.n12 dvss.t4 292.5
R1607 dvss.n11 dvss.t4 292.5
R1608 dvss.n26 dvss.n25 252.459
R1609 dvss.n6 dvss.t1 239.136
R1610 dvss.t2 dvss.n42 233.216
R1611 dvss.n1 dvss.t7 229.315
R1612 dvss.n34 dvss.n33 195.184
R1613 dvss.n66 dvss.n65 195
R1614 dvss.n65 dvss.n64 195
R1615 dvss.n37 dvss.n36 195
R1616 dvss.n38 dvss.n37 195
R1617 dvss.n35 dvss.n32 195
R1618 dvss.n43 dvss.n35 195
R1619 dvss.n52 dvss.n22 195
R1620 dvss.n48 dvss.n22 195
R1621 dvss.n28 dvss.n21 195
R1622 dvss.n23 dvss.n21 195
R1623 dvss.n23 dvss.n19 155.083
R1624 dvss.n24 dvss.n14 146.25
R1625 dvss.n25 dvss.n24 146.25
R1626 dvss.n62 dvss.n61 146.25
R1627 dvss.n63 dvss.n62 146.25
R1628 dvss.n61 dvss.n60 138.166
R1629 dvss.n53 dvss.n52 116.504
R1630 dvss.t0 dvss.t3 100.984
R1631 dvss.n47 dvss.n46 97.6305
R1632 dvss.n61 dvss.n13 86.5887
R1633 dvss.n36 dvss.n8 86.1306
R1634 dvss.n3 dvss.t5 84.1047
R1635 dvss.n39 dvss.n33 81.8974
R1636 dvss.n36 dvss.n7 74.9169
R1637 dvss.n45 dvss.n33 74.0493
R1638 dvss.n52 dvss.n51 57.0188
R1639 dvss.n58 dvss.n57 55.3148
R1640 dvss.n53 dvss.n29 53.0829
R1641 dvss.n60 dvss.n59 53.0829
R1642 dvss.n50 dvss.n47 48.155
R1643 dvss.n55 dvss.n19 46.8857
R1644 dvss.n39 dvss.n32 43.9756
R1645 dvss.n51 dvss.n50 42.7064
R1646 dvss.n66 dvss.n8 39.1038
R1647 dvss.n30 dvss.n16 31.8699
R1648 dvss.n57 dvss.n16 26.2862
R1649 dvss.n68 dvss.n67 17.1865
R1650 dvss.n46 dvss.n45 17.0668
R1651 dvss.n29 dvss.n6 14.0183
R1652 dvss.n68 dvss.n7 13.3694
R1653 dvss.n46 dvss.n32 12.1441
R1654 dvss.n27 dvss.n16 11.3033
R1655 dvss.n59 dvss.n58 10.109
R1656 dvss.n51 dvss.n31 6.79342
R1657 dvss.n59 dvss.n14 6.606
R1658 dvss.n5 dvss.n0 5.813
R1659 dvss.n58 dvss.n15 5.62852
R1660 dvss.n13 dvss.n2 5.6005
R1661 dvss.n29 dvss.n28 4.75646
R1662 dvss.n67 dvss.n1 4.6505
R1663 dvss.n67 dvss.n66 2.95435
R1664 dvss.n3 dvss.n0 2.6255
R1665 dvss.n70 dvss.n2 2.33934
R1666 dvss.n27 dvss.n2 1.88621
R1667 dvss.n69 dvss.n68 1.82171
R1668 dvss.n31 dvss.n30 1.46336
R1669 dvss.n69 dvss.n6 1.44933
R1670 dvss.n4 dvss.n3 1.2505
R1671 dvss.n47 dvss.n15 1.09622
R1672 dvss.n5 dvss 0.8755
R1673 dvss.n4 dvss 0.583833
R1674 dvss.n72 dvss.n0 0.438
R1675 dvss.n28 dvss.n27 0.26472
R1676 dvss.n69 dvss 0.119327
R1677 dvss.n70 dvss.n69 0.0769887
R1678 dvss.n16 dvss.n14 0.0592156
R1679 dvss.n71 dvss.n1 0.0536915
R1680 dvss.n70 dvss.n5 0.0472557
R1681 dvss.n71 dvss.n70 0.0133337
R1682 dvss.n72 dvss.n71 0.0125637
R1683 dvss.n5 dvss.n4 0.0019313
R1684 dvss dvss.n72 0.00178337
R1685 dvss.n4 dvss 0.000977099
R1686 dout.n1 dout.t0 243.876
R1687 dout.n0 dout.t1 230.631
R1688 dout.n0 dout.t2 228.215
R1689 dout.n1 dout.n0 3.11789
R1690 dout dout.n1 0.306432
R1691 a_2982_4700.t1 a_2982_4700.n0 661.461
R1692 a_2982_4700.n0 a_2982_4700.t0 236.12
R1693 a_2982_4700.n0 a_2982_4700.t3 108.308
R1694 a_2982_4700.n0 a_2982_4700.t5 107.8
R1695 a_2982_4700.n1 a_2982_4700.t2 107.362
R1696 a_2982_4700.n1 a_2982_4700.t4 105.01
R1697 a_2982_4700.n0 a_2982_4700.n1 16.7414
C0 a_866_518# a_534_518# 0.307869f
C1 a_5826_9768# a_5494_9768# 0.307869f
C2 a_10806_9768# a_11138_9768# 0.307869f
C3 rc_osc_level_shifter_0.out_h a_8714_4659# 0.326647f
C4 a_6676_3118# a_7008_3118# 0.307869f
C5 a_11304_7168# avdd 0.516263f
C6 a_11138_9768# a_11470_9768# 0.307869f
C7 dout a_7718_4786# 1.09434f
C8 rc_osc_level_shifter_0.outb_h a_7718_4786# 0.183562f
C9 a_5514_518# a_5846_518# 0.307869f
C10 a_4830_9768# avss 0.142763f
C11 a_4518_518# a_4850_518# 0.307869f
C12 a_7174_518# avss 0.184675f
C13 a_9996_3118# a_10328_3118# 0.307869f
C14 a_5660_7168# a_5328_7168# 0.307869f
C15 avdd a_3004_7168# 0.548273f
C16 avdd a_7718_4786# 0.60786f
C17 a_2526_518# a_2858_518# 0.307869f
C18 a_5826_9768# avss 0.142763f
C19 a_11636_7168# rc_osc_level_shifter_0.inb_l 0.164792f
C20 a_680_7168# a_1012_7168# 0.307869f
C21 a_5348_3118# a_5016_3118# 0.307869f
C22 a_8980_7168# avss 0.243852f
C23 a_9664_3118# avss 0.211499f
C24 a_3502_9768# a_3834_9768# 0.307869f
C25 a_6656_7168# a_6324_7168# 0.307869f
C26 ena a_7718_4786# 0.523822f
C27 avss a_10162_518# 0.184675f
C28 a_11636_7168# avss 0.808235f
C29 a_4000_7168# avdd 0.385508f
C30 a_7818_9768# avss 0.142763f
C31 a_5348_3118# avss 0.694407f
C32 a_11324_3118# avss 0.20921f
C33 a_10660_3118# avss 0.20921f
C34 a_6656_7168# avdd 0.548273f
C35 a_5846_518# a_6178_518# 0.307869f
C36 a_2672_7168# avdd 0.548273f
C37 a_6676_3118# avss 0.739782f
C38 a_8004_3118# avss 0.243263f
C39 a_3854_518# avss 0.184675f
C40 a_6158_9768# avss 0.142763f
C41 a_9830_518# avss 0.184675f
C42 rc_osc_level_shifter_0.out_h a_5862_4788# 0.164806f
C43 a_3336_7168# avdd 0.548273f
C44 a_8316_7168# a_8648_7168# 0.307869f
C45 a_10328_3118# avss 0.20921f
C46 a_7486_9768# avss 0.142763f
C47 a_5992_7168# a_6324_7168# 0.307869f
C48 a_5826_9768# a_6158_9768# 0.307869f
C49 a_6842_518# avss 0.184675f
C50 avdd a_10972_7168# 0.609955f
C51 a_3480_4788# avss 0.828006f
C52 a_8714_4659# rc_osc_level_shifter_0.outb_h 0.229072f
C53 a_11158_518# a_10826_518# 0.307869f
C54 a_11324_3118# a_11636_7168# 0.325625f
C55 a_3522_518# avss 0.184675f
C56 a_11304_7168# avss 0.145925f
C57 a_7174_518# a_6842_518# 0.307869f
C58 rc_osc_level_shifter_0.inb_l a_7718_4786# 0.881308f
C59 a_10806_9768# avss 0.142763f
C60 a_1344_7168# a_1012_7168# 0.307869f
C61 a_1862_518# avss 0.184675f
C62 a_5992_7168# avdd 0.548273f
C63 a_8714_4659# avdd 0.401456f
C64 a_11470_9768# avss 0.307678f
C65 avdd a_4352_3118# 0.307869f
C66 avdd a_2340_7168# 0.399783f
C67 a_2858_518# avss 0.184675f
C68 a_4996_7168# a_4664_7168# 0.307869f
C69 a_9830_518# a_10162_518# 0.307869f
C70 a_3004_7168# avss 0.209517f
C71 avss a_7718_4786# 0.630608f
C72 a_6656_7168# a_6988_7168# 0.307869f
C73 a_2526_4188# avss 0.699047f
C74 a_7154_9768# avss 0.142763f
C75 a_4996_7168# avss 0.209517f
C76 a_6012_3118# avss 0.739782f
C77 a_9332_3118# avss 0.214403f
C78 a_10640_7168# a_10972_7168# 0.307869f
C79 a_7486_9768# a_7818_9768# 0.307869f
C80 a_10660_3118# a_10328_3118# 0.307869f
C81 a_11304_7168# a_11636_7168# 0.307345f
C82 a_6260_4788# avss 0.892467f
C83 a_1842_9768# a_2174_9768# 0.307869f
C84 a_3190_518# avss 0.184675f
C85 a_8834_518# avss 0.184675f
C86 a_4000_7168# avss 0.209517f
C87 a_4854_5653# avdd 0.680997f
C88 a_4684_3118# a_4352_3118# 0.307869f
C89 a_6344_3118# avss 0.739782f
C90 a_6656_7168# avss 0.209517f
C91 a_8502_518# a_8170_518# 0.307869f
C92 a_5846_518# avss 0.184675f
C93 avdd a_5470_5653# 0.761298f
C94 a_5660_7168# avdd 0.548273f
C95 a_2672_7168# avss 0.209517f
C96 a_3502_9768# a_3170_9768# 0.307869f
C97 a_9478_9768# a_9810_9768# 0.307869f
C98 a_3854_518# a_3522_518# 0.307869f
C99 a_9664_3118# a_9332_3118# 0.307869f
C100 a_6490_9768# a_6822_9768# 0.307869f
C101 a_5862_4788# rc_osc_level_shifter_0.outb_h 0.140134f
C102 a_4186_518# avss 0.184675f
C103 a_1178_9768# a_846_9768# 0.307869f
C104 a_3336_7168# avss 0.209517f
C105 a_1510_9768# avss 0.142763f
C106 a_4592_4788# avss 0.824116f
C107 a_5862_4788# avdd 0.82569f
C108 a_4166_9768# a_3834_9768# 0.307869f
C109 avss a_10972_7168# 0.144844f
C110 a_2526_518# a_2194_518# 0.307869f
C111 a_7340_3118# a_7672_3118# 0.307869f
C112 a_1842_9768# avss 0.142763f
C113 a_10142_9768# a_9810_9768# 0.307869f
C114 a_1178_9768# avss 0.142763f
C115 a_5992_7168# avss 0.209517f
C116 a_7672_3118# avss 0.285635f
C117 a_5680_3118# avss 0.739782f
C118 a_2340_7168# avss 0.209517f
C119 avss a_4352_3118# 0.356069f
C120 a_7154_9768# a_7486_9768# 0.307869f
C121 a_3502_9768# avss 0.142763f
C122 a_8668_3118# avss 0.218069f
C123 a_8502_518# avss 0.184675f
C124 a_7652_7168# a_7320_7168# 0.307869f
C125 a_6988_7168# a_7320_7168# 0.307869f
C126 a_7652_7168# a_7984_7168# 0.307869f
C127 a_6344_3118# a_6676_3118# 0.307869f
C128 a_11158_518# avss 0.184675f
C129 a_5328_7168# avdd 0.436049f
C130 dout dvdd 0.892013f
C131 a_8336_3118# avss 0.221431f
C132 a_4850_518# a_5182_518# 0.307869f
C133 a_534_518# avss 0.348434f
C134 a_4186_518# a_3854_518# 0.307869f
C135 a_3522_518# a_3190_518# 0.307869f
C136 dvdd avdd 1.48803f
C137 a_1676_7168# a_2008_7168# 0.307869f
C138 avdd a_3668_7168# 0.548273f
C139 avss a_9810_9768# 0.142763f
C140 avss a_7320_7168# 0.209517f
C141 a_7984_7168# avss 0.209517f
C142 rc_osc_level_shifter_0.out_h rc_osc_level_shifter_0.outb_h 3.79716f
C143 avss a_1012_7168# 0.239502f
C144 a_3190_518# a_2858_518# 0.307869f
C145 a_5660_7168# avss 0.209517f
C146 a_9146_9768# a_8814_9768# 0.307869f
C147 a_5148_4788# avss 0.865328f
C148 a_5348_3118# a_5680_3118# 0.307869f
C149 rc_osc_level_shifter_0.out_h avdd 2.25409f
C150 dvdd ena 1.57004f
C151 a_5862_4788# a_6702_5653# 0.11184f
C152 a_4166_9768# a_4498_9768# 0.307869f
C153 a_8316_7168# avss 0.243852f
C154 a_8004_3118# a_7672_3118# 0.307869f
C155 a_2672_7168# a_3004_7168# 0.307869f
C156 a_4332_7168# a_4664_7168# 0.307869f
C157 a_5862_4788# avss 1.04053f
C158 a_4518_518# avss 0.184675f
C159 a_2194_518# avss 0.184675f
C160 a_1198_518# a_866_518# 0.307869f
C161 rc_osc_level_shifter_0.out_h ena 0.3516f
C162 a_10142_9768# a_10474_9768# 0.307869f
C163 a_6822_9768# avss 0.142763f
C164 a_3006_5653# avdd 0.816596f
C165 a_6344_3118# a_6012_3118# 0.307869f
C166 a_11304_7168# a_10972_7168# 0.307869f
C167 a_9166_518# a_9498_518# 0.307869f
C168 a_8482_9768# a_8150_9768# 0.307869f
C169 a_3336_7168# a_3004_7168# 0.307869f
C170 a_8004_3118# a_8336_3118# 0.307869f
C171 a_4332_7168# avss 0.209517f
C172 a_4850_518# avss 0.184675f
C173 a_2838_9768# a_3170_9768# 0.307869f
C174 a_846_9768# a_514_9768# 0.307869f
C175 a_9146_9768# a_9478_9768# 0.307869f
C176 a_10992_3118# avss 0.20921f
C177 a_9644_7168# a_9312_7168# 0.307869f
C178 a_1676_7168# a_1344_7168# 0.307869f
C179 a_9000_3118# avss 0.215228f
C180 a_5328_7168# avss 0.209517f
C181 dvdd rc_osc_level_shifter_0.inb_l 0.663728f
C182 a_514_9768# avss 0.305402f
C183 a_866_518# avss 0.184675f
C184 a_2506_9768# a_2838_9768# 0.307869f
C185 a_1198_518# a_1530_518# 0.307869f
C186 a_11490_518# avss 0.348069f
C187 a_8150_9768# avss 0.142763f
C188 avss a_10474_9768# 0.142763f
C189 a_6012_3118# a_5680_3118# 0.307869f
C190 a_10494_518# a_10826_518# 0.307869f
C191 dvdd avss 1.32652f
C192 a_680_7168# avss 0.238959f
C193 rc_osc_level_shifter_0.out_h rc_osc_level_shifter_0.inb_l 0.255743f
C194 a_3668_7168# avss 0.209517f
C195 a_2008_7168# avss 0.209517f
C196 a_2838_9768# avss 0.142763f
C197 a_6324_7168# avdd 0.548273f
C198 a_5514_518# a_5182_518# 0.307869f
C199 dout avdd 0.101166f
C200 a_11890_5939# dvdd 0.120615f
C201 a_9644_7168# avdd 0.305891f
C202 a_5704_4788# avss 0.86884f
C203 avdd rc_osc_level_shifter_0.outb_h 1.60324f
C204 a_8502_518# a_8834_518# 0.307869f
C205 rc_osc_level_shifter_0.out_h avss 4.2566f
C206 a_4166_9768# avss 0.142763f
C207 a_6510_518# a_6178_518# 0.307869f
C208 a_2672_7168# a_2340_7168# 0.307869f
C209 a_10992_3118# a_11324_3118# 0.307869f
C210 a_1510_9768# a_1842_9768# 0.307869f
C211 a_10992_3118# a_10660_3118# 0.307869f
C212 dout ena 0.18382f
C213 a_8648_7168# avss 0.243852f
C214 a_1178_9768# a_1510_9768# 0.307869f
C215 ena rc_osc_level_shifter_0.outb_h 0.463304f
C216 a_1530_518# avss 0.184675f
C217 a_8150_9768# a_7818_9768# 0.307869f
C218 a_8482_9768# a_8814_9768# 0.307869f
C219 dvdd a_11636_7168# 1.06568f
C220 a_1862_518# a_2194_518# 0.307869f
C221 ena avdd 1.6305f
C222 a_3834_9768# avss 0.142763f
C223 a_7560_4786# ena 0.161553f
C224 a_9146_9768# avss 0.142763f
C225 a_7838_518# a_8170_518# 0.307869f
C226 a_7506_518# a_7838_518# 0.307869f
C227 a_7154_9768# a_6822_9768# 0.307869f
C228 a_8980_7168# a_8648_7168# 0.307869f
C229 a_10640_7168# avdd 0.609955f
C230 a_9166_518# avss 0.184675f
C231 a_9482_5327# rc_osc_level_shifter_0.out_h 0.102468f
C232 a_5514_518# avss 0.184675f
C233 avss a_1344_7168# 0.239502f
C234 a_5862_4788# a_6260_4788# 0.175672f
C235 a_5494_9768# a_5162_9768# 0.307869f
C236 a_9312_7168# avss 0.243852f
C237 a_8814_9768# avss 0.142763f
C238 a_6988_7168# avdd 0.342919f
C239 dout rc_osc_level_shifter_0.inb_l 0.13931f
C240 a_10806_9768# a_10474_9768# 0.307869f
C241 a_8668_3118# a_8336_3118# 0.307869f
C242 a_4000_7168# a_4332_7168# 0.307869f
C243 rc_osc_level_shifter_0.inb_l rc_osc_level_shifter_0.outb_h 0.228327f
C244 a_9498_518# avss 0.184675f
C245 a_10308_7168# avdd 0.609955f
C246 a_10826_518# avss 0.184675f
C247 a_9644_7168# a_9976_7168# 0.307869f
C248 a_9000_3118# a_9332_3118# 0.307869f
C249 a_6324_7168# avss 0.209517f
C250 a_5162_9768# avss 0.142763f
C251 a_4996_7168# a_5328_7168# 0.307869f
C252 a_6490_9768# avss 0.142763f
C253 rc_osc_level_shifter_0.inb_l avdd 0.368358f
C254 avdd a_6702_5653# 0.791907f
C255 a_7838_518# avss 0.184675f
C256 a_4186_518# a_4518_518# 0.307869f
C257 a_9644_7168# avss 0.198487f
C258 a_2924_4788# avss 0.868706f
C259 rc_osc_level_shifter_0.outb_h avss 4.51566f
C260 a_4830_9768# a_5162_9768# 0.307869f
C261 dvdd a_7718_4786# 1.2174f
C262 avdd a_3622_5653# 0.790633f
C263 a_9976_7168# avdd 0.609955f
C264 a_8980_7168# a_9312_7168# 0.307869f
C265 a_5660_7168# a_5992_7168# 0.307869f
C266 a_6510_518# avss 0.184675f
C267 a_4036_4788# avss 0.823951f
C268 a_11138_9768# avss 0.142763f
C269 a_1676_7168# avss 0.228829f
C270 a_10494_518# avss 0.184675f
C271 a_11890_5939# dout 0.638473f
C272 a_6178_518# avss 0.184675f
C273 avdd avss 0.355979p
C274 a_7560_4786# avss 0.445517f
C275 ena rc_osc_level_shifter_0.inb_l 1.01705f
C276 avss a_4498_9768# 0.142763f
C277 a_2526_518# avss 0.184675f
C278 rc_osc_level_shifter_0.out_h a_7718_4786# 0.144107f
C279 rc_osc_level_shifter_0.out_h a_2526_4188# 0.106807f
C280 a_9478_9768# avss 0.142763f
C281 a_4830_9768# a_4498_9768# 0.307869f
C282 a_1862_518# a_1530_518# 0.307869f
C283 a_10640_7168# a_10308_7168# 0.307869f
C284 ena avss 1.15253f
C285 a_4000_7168# a_3668_7168# 0.307869f
C286 a_7340_3118# a_7008_3118# 0.307869f
C287 a_5016_3118# a_4684_3118# 0.307869f
C288 a_9996_3118# avss 0.20921f
C289 a_6086_5653# avdd 0.788381f
C290 a_2506_9768# a_2174_9768# 0.307869f
C291 a_11890_5939# ena 0.177772f
C292 a_5182_518# avss 0.184675f
C293 a_7008_3118# avss 0.550938f
C294 a_10494_518# a_10162_518# 0.307869f
C295 a_10640_7168# avss 0.144844f
C296 a_4684_3118# avss 0.339621f
C297 a_11636_7168# avdd 1.3903f
C298 a_9482_5327# rc_osc_level_shifter_0.outb_h 0.202516f
C299 avss a_8170_518# 0.184675f
C300 a_9498_518# a_9830_518# 0.307869f
C301 a_7506_518# avss 0.184675f
C302 a_10142_9768# avss 0.142763f
C303 avss a_3170_9768# 0.142763f
C304 a_8316_7168# a_7984_7168# 0.307869f
C305 a_2174_9768# avss 0.142763f
C306 a_6490_9768# a_6158_9768# 0.307869f
C307 a_3336_7168# a_3668_7168# 0.307869f
C308 a_1198_518# avss 0.184675f
C309 a_8482_9768# avss 0.142763f
C310 a_9482_5327# avdd 0.528099f
C311 a_7506_518# a_7174_518# 0.307869f
C312 a_8668_3118# a_9000_3118# 0.307869f
C313 a_9996_3118# a_9664_3118# 0.307869f
C314 a_7652_7168# avss 0.209517f
C315 a_6988_7168# avss 0.209517f
C316 a_10308_7168# a_9976_7168# 0.307869f
C317 a_846_9768# avss 0.142763f
C318 a_10308_7168# avss 0.144844f
C319 a_5494_9768# avss 0.142763f
C320 a_9482_5327# ena 0.117123f
C321 a_5016_3118# avss 0.401051f
C322 rc_osc_level_shifter_0.inb_l avss 0.875565f
C323 a_6510_518# a_6842_518# 0.307869f
C324 a_11490_518# a_11158_518# 0.307869f
C325 a_2506_9768# avss 0.142763f
C326 a_7340_3118# avss 0.349196f
C327 a_4664_7168# avss 0.209517f
C328 a_2008_7168# a_2340_7168# 0.307869f
C329 a_4238_5653# avdd 0.701946f
C330 a_9166_518# a_8834_518# 0.307869f
C331 a_9976_7168# avss 0.144844f
C332 dout dvss 1.18563f
C333 ena dvss 1.822f
C334 dvdd dvss 6.22115f
C335 avss dvss 6.804884f
C336 avdd dvss 0.394817p
C337 a_11490_518# dvss 0.297186f
C338 a_11324_3118# dvss 0.241933f
C339 a_11158_518# dvss 0.261223f
C340 a_10992_3118# dvss 0.241933f
C341 a_10826_518# dvss 0.261223f
C342 a_10660_3118# dvss 0.241933f
C343 a_10494_518# dvss 0.261223f
C344 a_10328_3118# dvss 0.254752f
C345 a_10162_518# dvss 0.261223f
C346 a_9996_3118# dvss 0.255929f
C347 a_9830_518# dvss 0.261223f
C348 a_9664_3118# dvss 0.241933f
C349 a_9498_518# dvss 0.261223f
C350 a_9332_3118# dvss 0.241933f
C351 a_9166_518# dvss 0.261223f
C352 a_9000_3118# dvss 0.241933f
C353 a_8834_518# dvss 0.261223f
C354 a_8668_3118# dvss 0.241933f
C355 a_8502_518# dvss 0.261223f
C356 a_8336_3118# dvss 0.241933f
C357 a_8170_518# dvss 0.261223f
C358 a_8004_3118# dvss 0.241933f
C359 a_7838_518# dvss 0.261223f
C360 a_7672_3118# dvss 0.241933f
C361 a_7506_518# dvss 0.261223f
C362 a_7340_3118# dvss 0.241933f
C363 a_7174_518# dvss 0.261223f
C364 a_7008_3118# dvss 0.241933f
C365 a_6842_518# dvss 0.261223f
C366 a_6676_3118# dvss 0.241933f
C367 a_6510_518# dvss 0.261223f
C368 a_6344_3118# dvss 0.241933f
C369 a_6178_518# dvss 0.261223f
C370 a_6012_3118# dvss 0.241933f
C371 a_5846_518# dvss 0.261223f
C372 a_5680_3118# dvss 0.241933f
C373 a_5514_518# dvss 0.261223f
C374 a_5348_3118# dvss 0.241933f
C375 a_5182_518# dvss 0.261223f
C376 a_5016_3118# dvss 0.241933f
C377 a_4850_518# dvss 0.261223f
C378 a_4684_3118# dvss 0.241933f
C379 a_4518_518# dvss 0.261223f
C380 a_4352_3118# dvss 0.241933f
C381 a_4186_518# dvss 0.261223f
C382 a_3854_518# dvss 0.261223f
C383 a_3522_518# dvss 0.261223f
C384 a_3190_518# dvss 0.261223f
C385 a_2858_518# dvss 0.261223f
C386 a_2526_518# dvss 0.261223f
C387 a_2194_518# dvss 0.261223f
C388 a_1862_518# dvss 0.261223f
C389 a_1530_518# dvss 0.261223f
C390 a_1198_518# dvss 0.261223f
C391 a_866_518# dvss 0.261223f
C392 a_534_518# dvss 0.296272f
C393 a_11890_5939# dvss 0.633389f
C394 rc_osc_level_shifter_0.outb_h dvss 5.057272f
C395 rc_osc_level_shifter_0.inb_l dvss 0.970466f
C396 a_7718_4786# dvss 0.857037f
C397 a_5862_4788# dvss 0.146786f
C398 rc_osc_level_shifter_0.out_h dvss 5.442275f
C399 a_11636_7168# dvss 2.90914f
C400 a_11470_9768# dvss 0.296245f
C401 a_11304_7168# dvss 0.241107f
C402 a_11138_9768# dvss 0.261295f
C403 a_10972_7168# dvss 0.240839f
C404 a_10806_9768# dvss 0.261295f
C405 a_10640_7168# dvss 0.240839f
C406 a_10474_9768# dvss 0.261295f
C407 a_10308_7168# dvss 0.240839f
C408 a_10142_9768# dvss 0.261295f
C409 a_9976_7168# dvss 0.240839f
C410 a_9810_9768# dvss 0.261295f
C411 a_9644_7168# dvss 0.242958f
C412 a_9478_9768# dvss 0.261295f
C413 a_9312_7168# dvss 0.240839f
C414 a_9146_9768# dvss 0.261295f
C415 a_8980_7168# dvss 0.240839f
C416 a_8814_9768# dvss 0.261295f
C417 a_8648_7168# dvss 0.240839f
C418 a_8482_9768# dvss 0.261295f
C419 a_8316_7168# dvss 0.240839f
C420 a_8150_9768# dvss 0.261295f
C421 a_7984_7168# dvss 0.240839f
C422 a_7818_9768# dvss 0.261295f
C423 a_7652_7168# dvss 0.240839f
C424 a_7486_9768# dvss 0.261295f
C425 a_7320_7168# dvss 0.240839f
C426 a_7154_9768# dvss 0.261295f
C427 a_6988_7168# dvss 0.240839f
C428 a_6822_9768# dvss 0.261295f
C429 a_6656_7168# dvss 0.240839f
C430 a_6490_9768# dvss 0.261295f
C431 a_6324_7168# dvss 0.240839f
C432 a_6158_9768# dvss 0.261295f
C433 a_5992_7168# dvss 0.240839f
C434 a_5826_9768# dvss 0.261295f
C435 a_5660_7168# dvss 0.240839f
C436 a_5494_9768# dvss 0.261295f
C437 a_5328_7168# dvss 0.240839f
C438 a_5162_9768# dvss 0.261295f
C439 a_4996_7168# dvss 0.240839f
C440 a_4830_9768# dvss 0.261295f
C441 a_4664_7168# dvss 0.240839f
C442 a_4498_9768# dvss 0.261295f
C443 a_4332_7168# dvss 0.240839f
C444 a_4166_9768# dvss 0.261295f
C445 a_4000_7168# dvss 0.240839f
C446 a_3834_9768# dvss 0.261295f
C447 a_3668_7168# dvss 0.240839f
C448 a_3502_9768# dvss 0.261295f
C449 a_3336_7168# dvss 0.240839f
C450 a_3170_9768# dvss 0.261295f
C451 a_3004_7168# dvss 0.240839f
C452 a_2838_9768# dvss 0.261295f
C453 a_2672_7168# dvss 0.240839f
C454 a_2506_9768# dvss 0.261295f
C455 a_2340_7168# dvss 0.240839f
C456 a_2174_9768# dvss 0.261295f
C457 a_2008_7168# dvss 0.240839f
C458 a_1842_9768# dvss 0.261295f
C459 a_1676_7168# dvss 0.240839f
C460 a_1510_9768# dvss 0.261295f
C461 a_1344_7168# dvss 0.240839f
C462 a_1178_9768# dvss 0.261295f
C463 a_1012_7168# dvss 0.240839f
C464 a_846_9768# dvss 0.261295f
C465 a_680_7168# dvss 0.240839f
C466 a_514_9768# dvss 0.297362f
C467 a_2982_4700.n0 dvss 2.14348f
C468 a_2982_4700.t3 dvss 0.165851f
C469 a_2982_4700.t5 dvss 0.164149f
C470 a_2982_4700.t2 dvss 0.162716f
C471 a_2982_4700.t4 dvss 0.153424f
C472 a_2982_4700.n1 dvss 1.14864f
C473 a_5306_4788.t2 dvss 3.67495f
C474 a_514_7168.t1 dvss 2.3123f
C475 a_1414_4786.n0 dvss 7.603701f
C476 a_1414_4786.t4 dvss 0.349517f
C477 a_1414_4786.t6 dvss 0.342485f
C478 a_1414_4786.t5 dvss 0.342485f
C479 a_1414_4786.t8 dvss 0.342485f
C480 a_1414_4786.t11 dvss 0.342485f
C481 a_1414_4786.t7 dvss 0.342485f
C482 a_1414_4786.t10 dvss 0.342485f
C483 a_1414_4786.t9 dvss 0.342485f
C484 a_1414_4786.t1 dvss 0.342485f
C485 a_4750_4788.t2 dvss 3.67205f
C486 rc_osc_level_shifter_0.out_h.n0 dvss 3.99803f
C487 rc_osc_level_shifter_0.out_h.t5 dvss 0.266754f
C488 rc_osc_level_shifter_0.out_h.t4 dvss 0.310921f
C489 rc_osc_level_shifter_0.out_h.t6 dvss 0.259169f
C490 rc_osc_level_shifter_0.out_h.t3 dvss 0.252779f
C491 rc_osc_level_shifter_0.out_h.t2 dvss 0.283777f
C492 a_3082_4788.t2 dvss 3.38418f
C493 rc_osc_level_shifter_0.outb_h.n0 dvss 2.27957f
C494 rc_osc_level_shifter_0.outb_h.t2 dvss 0.661159f
C495 rc_osc_level_shifter_0.outb_h.t3 dvss 0.315276f
C496 rc_osc_level_shifter_0.outb_h.t4 dvss 0.273065f
C497 a_2368_4788.n0 dvss 4.61781f
C498 a_2368_4788.n1 dvss 1.89182f
C499 a_2368_4788.t2 dvss 0.32443f
C500 a_2368_4788.t7 dvss 0.32443f
C501 a_2368_4788.t6 dvss 0.32443f
C502 a_2368_4788.t8 dvss 0.32443f
C503 a_2368_4788.t4 dvss 0.32443f
C504 a_2368_4788.t5 dvss 0.32443f
C505 a_2368_4788.t10 dvss 0.32443f
C506 a_2368_4788.t9 dvss 0.331908f
C507 a_4194_4788.t3 dvss 3.57171f
C508 a_3638_4788.t3 dvss 3.57318f
C509 avdd.n0 dvss 0.977171f
C510 avdd.n1 dvss 0.534269f
C511 avdd.n2 dvss 0.534269f
C512 avdd.n3 dvss 0.534269f
C513 avdd.n4 dvss 0.534269f
C514 avdd.n5 dvss 0.534269f
C515 avdd.n6 dvss 0.534269f
C516 avdd.n7 dvss 0.534269f
C517 avdd.n8 dvss 0.534269f
C518 avdd.n9 dvss 0.534269f
C519 avdd.n10 dvss 0.534269f
C520 avdd.n11 dvss 0.534269f
C521 avdd.n12 dvss 0.534269f
C522 avdd.n13 dvss 0.534269f
C523 avdd.n14 dvss 0.534269f
C524 avdd.n15 dvss 0.534269f
C525 avdd.n16 dvss 0.534269f
C526 avdd.n17 dvss 0.534269f
C527 avdd.n18 dvss 0.534269f
C528 avdd.n19 dvss 0.534269f
C529 avdd.n20 dvss 0.534269f
C530 avdd.n21 dvss 2.62257f
C531 avdd.n22 dvss 9.08475f
C532 avdd.n23 dvss 6.14943f
C533 avdd.n24 dvss 3.96681f
C534 avdd.n25 dvss 0.637662f
C535 avdd.n26 dvss 0.433226f
C536 avdd.n27 dvss 0.433226f
C537 avdd.n29 dvss 0.127141f
C538 avdd.n32 dvss 0.127141f
C539 avdd.n33 dvss 0.116184f
C540 avdd.n34 dvss 0.116115f
C541 avdd.n35 dvss 0.116115f
C542 avdd.n36 dvss 1.19732f
C543 avdd.n37 dvss 0.116184f
C544 avdd.n38 dvss 1.19732f
C545 avdd.n39 dvss 0.116115f
C546 avdd.n40 dvss 0.116115f
C547 avdd.n41 dvss 0.15678f
C548 avdd.n42 dvss 0.15678f
C549 avdd.n43 dvss 0.116115f
C550 avdd.n44 dvss 0.116115f
C551 avdd.n45 dvss 1.19732f
C552 avdd.n46 dvss 0.116184f
C553 avdd.n47 dvss 0.116184f
C554 avdd.n48 dvss 1.19732f
C555 avdd.n50 dvss 0.116115f
C556 avdd.n53 dvss 0.108902f
C557 avdd.n54 dvss 0.116115f
C558 avdd.n58 dvss 0.245713f
C559 avdd.n59 dvss 0.116115f
C560 avdd.n60 dvss 0.116115f
C561 avdd.n61 dvss 1.95195f
C562 avdd.n62 dvss 0.116184f
C563 avdd.n63 dvss 1.19732f
C564 avdd.n64 dvss 0.116184f
C565 avdd.n65 dvss 0.116115f
C566 avdd.n66 dvss 0.116115f
C567 avdd.n67 dvss 0.494773f
C568 avdd.n69 dvss 1.10514f
C569 avdd.n70 dvss 1.07554f
C570 avdd.n71 dvss 0.116115f
C571 avdd.n72 dvss 0.313288f
C572 avdd.n73 dvss 0.245713f
C573 avdd.n74 dvss 0.272286f
C574 avdd.n75 dvss 0.116184f
C575 avdd.n77 dvss 1.94968f
C576 avdd.t32 dvss 1.502f
C577 avdd.n78 dvss 0.116184f
C578 avdd.n79 dvss 0.129461f
C579 avdd.n80 dvss 0.334904f
C580 avdd.n82 dvss 0.335851f
C581 avdd.n84 dvss 0.127141f
C582 avdd.n85 dvss 0.108902f
C583 avdd.n87 dvss 0.210051f
C584 avdd.n88 dvss 0.225752f
C585 avdd.n90 dvss 0.15678f
C586 avdd.n91 dvss 0.148401f
C587 avdd.n92 dvss 0.116184f
C588 avdd.t23 dvss 1.26565f
C589 avdd.n93 dvss 0.116184f
C590 avdd.n94 dvss 0.148401f
C591 avdd.n95 dvss 0.157227f
C592 avdd.n96 dvss 0.157227f
C593 avdd.n97 dvss 0.148401f
C594 avdd.n98 dvss 0.157227f
C595 avdd.n99 dvss 0.157227f
C596 avdd.n100 dvss 0.148401f
C597 avdd.n101 dvss 0.157227f
C598 avdd.n102 dvss 0.157227f
C599 avdd.n103 dvss 0.116184f
C600 avdd.n104 dvss 0.116184f
C601 avdd.t5 dvss 1.26565f
C602 avdd.n105 dvss 0.116184f
C603 avdd.n107 dvss 0.116115f
C604 avdd.n108 dvss 0.116115f
C605 avdd.t12 dvss 1.26565f
C606 avdd.n109 dvss 0.116184f
C607 avdd.n110 dvss 0.116184f
C608 avdd.n111 dvss 0.129607f
C609 avdd.n112 dvss 1.51361f
C610 avdd.n113 dvss 0.101373f
C611 avdd.n114 dvss 0.15678f
C612 avdd.n115 dvss 0.15678f
C613 avdd.n116 dvss 0.433226f
C614 avdd.n117 dvss 0.127141f
C615 avdd.n118 dvss 0.148401f
C616 avdd.n120 dvss 0.157227f
C617 avdd.n121 dvss 0.116184f
C618 avdd.n123 dvss 1.19732f
C619 avdd.n124 dvss 0.148401f
C620 avdd.n125 dvss 0.15678f
C621 avdd.n126 dvss 0.108902f
C622 avdd.n128 dvss 0.433226f
C623 avdd.n129 dvss 0.108902f
C624 avdd.n130 dvss 0.157227f
C625 avdd.n131 dvss 0.116184f
C626 avdd.n132 dvss 0.116115f
C627 avdd.n133 dvss 0.148401f
C628 avdd.n134 dvss 1.19732f
C629 avdd.n135 dvss 0.116184f
C630 avdd.n136 dvss 0.116115f
C631 avdd.n137 dvss 0.116115f
C632 avdd.n138 dvss 0.15678f
C633 avdd.n141 dvss 0.15678f
C634 avdd.n142 dvss 0.116115f
C635 avdd.n143 dvss 0.116115f
C636 avdd.n144 dvss 1.19732f
C637 avdd.n145 dvss 0.116184f
C638 avdd.n146 dvss 0.116184f
C639 avdd.n147 dvss 1.19732f
C640 avdd.n148 dvss 0.127141f
C641 avdd.n150 dvss 0.116115f
C642 avdd.n153 dvss 0.127141f
C643 avdd.n154 dvss 0.687512f
C644 avdd.n155 dvss 2.44157f
C645 avdd.n156 dvss 0.116115f
C646 avdd.n159 dvss 0.25456f
C647 avdd.n160 dvss 0.116115f
C648 avdd.n161 dvss 0.116115f
C649 avdd.n162 dvss 1.19732f
C650 avdd.n163 dvss 0.116184f
C651 avdd.n164 dvss 1.19732f
C652 avdd.n165 dvss 0.116184f
C653 avdd.n166 dvss 0.116115f
C654 avdd.n167 dvss 0.116115f
C655 avdd.n168 dvss 0.15678f
C656 avdd.n169 dvss 0.115751f
C657 avdd.n171 dvss 0.130882f
C658 avdd.n172 dvss 0.277653f
C659 avdd.n174 dvss 0.25203f
C660 avdd.n175 dvss 0.243896f
C661 avdd.n176 dvss 0.116184f
C662 avdd.t0 dvss 1.26565f
C663 avdd.n177 dvss 0.116184f
C664 avdd.n178 dvss 0.245621f
C665 avdd.n179 dvss 0.157227f
C666 avdd.n180 dvss 0.157227f
C667 avdd.n181 dvss 0.148401f
C668 avdd.n182 dvss 0.157227f
C669 avdd.n183 dvss 0.157227f
C670 avdd.n185 dvss 0.225752f
C671 avdd.n186 dvss 0.210051f
C672 avdd.n187 dvss 0.433226f
C673 avdd.n188 dvss 1.1334f
C674 avdd.n189 dvss 0.58202f
C675 avdd.n190 dvss 0.210051f
C676 avdd.n191 dvss 0.225752f
C677 avdd.n192 dvss 0.108902f
C678 avdd.n193 dvss 0.116184f
C679 avdd.t4 dvss 1.26565f
C680 avdd.n194 dvss 0.116184f
C681 avdd.n195 dvss 0.148401f
C682 avdd.n196 dvss 0.15678f
C683 avdd.n197 dvss 0.15678f
C684 avdd.n198 dvss 0.148401f
C685 avdd.n199 dvss 0.116184f
C686 avdd.t15 dvss 1.26565f
C687 avdd.n200 dvss 0.116184f
C688 avdd.n201 dvss 0.116115f
C689 avdd.n203 dvss 0.127141f
C690 avdd.n204 dvss 0.210051f
C691 avdd.n205 dvss 0.225752f
C692 avdd.n207 dvss 0.116115f
C693 avdd.n208 dvss 1.19732f
C694 avdd.n209 dvss 0.116115f
C695 avdd.n210 dvss 0.116184f
C696 avdd.n211 dvss 0.148401f
C697 avdd.n212 dvss 0.157227f
C698 avdd.n213 dvss 0.157227f
C699 avdd.n215 dvss 0.225752f
C700 avdd.n216 dvss 0.210051f
C701 avdd.n218 dvss 0.116115f
C702 avdd.n219 dvss 1.19732f
C703 avdd.n220 dvss 1.19732f
C704 avdd.n221 dvss 0.116115f
C705 avdd.n222 dvss 0.116184f
C706 avdd.n223 dvss 0.116115f
C707 avdd.n224 dvss 1.19732f
C708 avdd.n225 dvss 0.116115f
C709 avdd.n227 dvss 0.127141f
C710 avdd.n228 dvss 0.433226f
C711 avdd.n229 dvss 0.210051f
C712 avdd.n230 dvss 0.225752f
C713 avdd.n231 dvss 0.108902f
C714 avdd.n232 dvss 0.116184f
C715 avdd.t38 dvss 1.26565f
C716 avdd.n233 dvss 0.116184f
C717 avdd.n234 dvss 0.148401f
C718 avdd.n235 dvss 0.15678f
C719 avdd.n236 dvss 0.15678f
C720 avdd.n237 dvss 0.148401f
C721 avdd.n238 dvss 0.116184f
C722 avdd.t37 dvss 1.26565f
C723 avdd.n239 dvss 0.116184f
C724 avdd.n240 dvss 0.108902f
C725 avdd.n241 dvss 0.225752f
C726 avdd.n242 dvss 0.210051f
C727 avdd.n243 dvss 0.433226f
C728 avdd.n244 dvss 1.1334f
C729 avdd.n245 dvss 2.70052f
C730 avdd.n246 dvss 5.38473f
C731 avdd.n247 dvss 2.74627f
C732 avdd.n248 dvss 5.92469f
C733 avdd.n249 dvss 1.0739f
C734 avdd.n250 dvss 3.10845f
C735 avdd.n251 dvss 0.891503f
C736 avdd.n252 dvss 13.325f
C737 avdd.n253 dvss 2.93304f
C738 avdd.n254 dvss 1.61179f
C739 avdd.n255 dvss 0.732695f
C740 avdd.n256 dvss 0.116184f
C741 avdd.n257 dvss 0.116184f
C742 avdd.n258 dvss 0.305123f
C743 avdd.n259 dvss 0.12963f
C744 avdd.n260 dvss 0.967933f
C745 avdd.n261 dvss 2.45157f
C746 avdd.n262 dvss 3.10861f
C747 avdd.n263 dvss 5.73656f
C748 avdd.n264 dvss 4.41051f
C749 avdd.n265 dvss 3.15478f
C750 avdd.n266 dvss 3.65309f
C751 avdd.n267 dvss 15.7673f
C752 avdd.n268 dvss 13.3258f
C753 avdd.n269 dvss 7.601171f
C754 avdd.n270 dvss 1.7736f
C755 avdd.n271 dvss 0.891342f
C756 avdd.n272 dvss 1.4813f
C757 avdd.n273 dvss 0.843118f
C758 avdd.n274 dvss 0.726483f
C759 avdd.n275 dvss 1.31759f
C760 avdd.n276 dvss 0.25477f
C761 avdd.n277 dvss 0.122298f
C762 avdd.n278 dvss 0.232632f
C763 avdd.n279 dvss 0.116115f
C764 avdd.n280 dvss 0.116115f
C765 avdd.n281 dvss 1.36563f
C766 avdd.n282 dvss 0.116184f
C767 avdd.n283 dvss 0.116184f
C768 avdd.n284 dvss 1.38627f
C769 avdd.n285 dvss 0.559697f
C770 avdd.n286 dvss 0.17729f
C771 avdd.n287 dvss 0.116184f
C772 avdd.n288 dvss 0.212288f
C773 avdd.n289 dvss 0.116115f
C774 avdd.n290 dvss 0.121908f
C775 avdd.n292 dvss 0.116184f
C776 avdd.t25 dvss 0.732695f
C777 avdd.t17 dvss 0.732695f
C778 avdd.n293 dvss 0.140855f
C779 avdd.n294 dvss 0.239503f
C780 avdd.n295 dvss 0.116115f
C781 avdd.n296 dvss 0.732695f
C782 avdd.n297 dvss 0.653577f
C783 avdd.n298 dvss 0.116115f
C784 avdd.n299 dvss 0.108902f
C785 avdd.n300 dvss 0.116115f
C786 avdd.n301 dvss 0.133261f
C787 avdd.n302 dvss 0.27665f
C788 avdd.n303 dvss 0.17501f
C789 avdd.n304 dvss 0.116115f
C790 avdd.n305 dvss 0.205765f
C791 avdd.n306 dvss 0.303752f
C792 avdd.n307 dvss 0.211546f
C793 avdd.n308 dvss 0.116184f
C794 avdd.t27 dvss 1.45999f
C795 avdd.n309 dvss 0.116184f
C796 avdd.n310 dvss 0.132753f
C797 avdd.n311 dvss 0.155919f
C798 avdd.n313 dvss -2.09062f
C799 avdd.n314 dvss 1.64106f
C800 avdd.n315 dvss 0.157974f
C801 avdd.n316 dvss 0.125651f
C802 avdd.n317 dvss 0.116115f
C803 avdd.n318 dvss 0.976926f
C804 avdd.n319 dvss 3.90698f
C805 avdd.n320 dvss 3.64356f
C806 avdd.n321 dvss 7.603859f
C807 avdd.n322 dvss 1.77424f
C808 avdd.n323 dvss 0.624266f
C809 avdd.n324 dvss 2.31105f
C810 avdd.n325 dvss 7.10226f
C811 avdd.n326 dvss 30.8011f
C812 avdd.n327 dvss 35.673702f
C813 avdd.n328 dvss 29.6884f
C814 avdd.n329 dvss 15.4209f
C815 avss.n0 dvss 6.29454f
C816 avss.n1 dvss 1.3779f
C817 avss.n2 dvss 1.97943f
C818 avss.n3 dvss 0.595594f
C819 avss.n4 dvss 0.595594f
C820 avss.t44 dvss 0.631727f
C821 avss.n7 dvss 0.149265f
C822 avss.n9 dvss 0.238581f
C823 avss.n10 dvss 0.140759f
C824 avss.n11 dvss 2.03759f
C825 avss.n12 dvss 10.448501f
C826 avss.n19 dvss 0.178308f
C827 avss.t91 dvss 1.2815f
C828 avss.t18 dvss 1.13711f
C829 avss.t108 dvss 1.14313f
C830 avss.n27 dvss 0.926533f
C831 avss.t94 dvss 1.27453f
C832 avss.n28 dvss 0.595594f
C833 avss.n29 dvss 0.595594f
C834 avss.n30 dvss 1.97795f
C835 avss.n31 dvss 1.89525f
C836 avss.n32 dvss 0.368279f
C837 avss.n33 dvss 0.205615f
C838 avss.n34 dvss 0.312475f
C839 avss.n35 dvss 0.406374f
C840 avss.n36 dvss 1.94186f
C841 avss.t107 dvss 1.37729f
C842 avss.t157 dvss 1.361f
C843 avss.t116 dvss 1.361f
C844 avss.t29 dvss 1.361f
C845 avss.t124 dvss 1.361f
C846 avss.t165 dvss 1.361f
C847 avss.t51 dvss 1.361f
C848 avss.t123 dvss 1.361f
C849 avss.t48 dvss 1.361f
C850 avss.t26 dvss 1.361f
C851 avss.t13 dvss 1.361f
C852 avss.t62 dvss 1.36293f
C853 avss.t65 dvss 1.46556f
C854 avss.t68 dvss 1.46377f
C855 avss.t87 dvss 1.46377f
C856 avss.t15 dvss 1.46377f
C857 avss.t159 dvss 1.33591f
C858 avss.t164 dvss 1.46417f
C859 avss.t11 dvss 1.46417f
C860 avss.t110 dvss 1.46417f
C861 avss.t98 dvss 1.46417f
C862 avss.t84 dvss 1.46417f
C863 avss.t7 dvss 1.46417f
C864 avss.t115 dvss 1.46417f
C865 avss.t137 dvss 1.46417f
C866 avss.t106 dvss 1.46417f
C867 avss.t69 dvss 1.46417f
C868 avss.t135 dvss 1.46417f
C869 avss.t128 dvss 1.46417f
C870 avss.t142 dvss 1.46417f
C871 avss.t140 dvss 1.46417f
C872 avss.t8 dvss 1.46417f
C873 avss.t150 dvss 1.46417f
C874 avss.t56 dvss 1.46417f
C875 avss.t99 dvss 1.46417f
C876 avss.t105 dvss 1.46417f
C877 avss.t49 dvss 1.46417f
C878 avss.t151 dvss 1.46417f
C879 avss.t53 dvss 1.46417f
C880 avss.t147 dvss 1.46417f
C881 avss.t54 dvss 1.46417f
C882 avss.t47 dvss 1.46417f
C883 avss.t36 dvss 1.46417f
C884 avss.t83 dvss 1.46417f
C885 avss.t60 dvss 1.09813f
C886 avss.n37 dvss 0.732085f
C887 avss.t153 dvss 1.09813f
C888 avss.t113 dvss 1.46417f
C889 avss.t12 dvss 1.46417f
C890 avss.t138 dvss 1.46417f
C891 avss.t35 dvss 1.46417f
C892 avss.t102 dvss 1.46418f
C893 avss.t127 dvss 1.46379f
C894 avss.t143 dvss 1.46377f
C895 avss.t34 dvss 1.46377f
C896 avss.t46 dvss 1.46377f
C897 avss.t125 dvss 1.46377f
C898 avss.t19 dvss 1.46377f
C899 avss.t64 dvss 1.46377f
C900 avss.t149 dvss 1.46377f
C901 avss.t129 dvss 1.46377f
C902 avss.t82 dvss 1.46377f
C903 avss.t93 dvss 0.859745f
C904 avss.n38 dvss 0.987216f
C905 avss.n43 dvss 0.156942f
C906 avss.n44 dvss 0.555193f
C907 avss.n46 dvss 0.922315f
C908 avss.n47 dvss 0.106821f
C909 avss.t41 dvss 0.320065f
C910 avss.t90 dvss 1.67483f
C911 avss.t14 dvss 1.04686f
C912 avss.n51 dvss 0.135654f
C913 avss.n53 dvss 0.541789f
C914 avss.t10 dvss 1.23337f
C915 avss.t132 dvss 1.21532f
C916 avss.n60 dvss 0.791852f
C917 avss.n64 dvss 0.414904f
C918 avss.n65 dvss 0.679424f
C919 avss.t146 dvss 1.2815f
C920 avss.t31 dvss 1.23337f
C921 avss.t163 dvss 1.11304f
C922 avss.t39 dvss 1.2815f
C923 avss.n87 dvss 0.177516f
C924 avss.n88 dvss 0.291278f
C925 avss.n89 dvss 0.314482f
C926 avss.t30 dvss 1.2815f
C927 avss.t109 dvss 1.18524f
C928 avss.t52 dvss 1.16117f
C929 avss.t145 dvss 1.2815f
C930 avss.t131 dvss 1.09499f
C931 avss.t104 dvss 1.11906f
C932 avss.n115 dvss 0.902467f
C933 avss.n116 dvss 0.878402f
C934 avss.t79 dvss 1.2815f
C935 avss.t126 dvss 1.2815f
C936 avss.t40 dvss 1.04686f
C937 avss.t67 dvss 1.16719f
C938 avss.n127 dvss 0.950599f
C939 avss.n128 dvss 0.83027f
C940 avss.t112 dvss 1.2815f
C941 avss.t71 dvss 1.2815f
C942 avss.n138 dvss 0.998731f
C943 avss.t33 dvss 0.782138f
C944 avss.n139 dvss 0.998731f
C945 avss.t28 dvss 1.2815f
C946 avss.t114 dvss 1.06491f
C947 avss.t76 dvss 0.998731f
C948 avss.n145 dvss 0.124635f
C949 avss.n146 dvss 0.132792f
C950 avss.n147 dvss 0.215298f
C951 avss.n148 dvss 0.21538f
C952 avss.n153 dvss 0.998731f
C953 avss.t89 dvss 0.631727f
C954 avss.n154 dvss 0.649777f
C955 avss.n155 dvss 0.499365f
C956 avss.t72 dvss 0.998731f
C957 avss.n171 dvss 2.69592f
C958 avss.n172 dvss 0.80824f
C959 avss.n176 dvss 0.998731f
C960 avss.t144 dvss 0.782138f
C961 avss.n177 dvss 0.998731f
C962 avss.n180 dvss 0.998731f
C963 avss.t96 dvss 0.782138f
C964 avss.n181 dvss 0.998731f
C965 avss.t1 dvss 0.998731f
C966 avss.n204 dvss 0.30263f
C967 avss.n210 dvss 0.998731f
C968 avss.t156 dvss 0.782138f
C969 avss.t59 dvss 1.2815f
C970 avss.n218 dvss 0.998731f
C971 avss.t50 dvss 0.782138f
C972 avss.n219 dvss 0.998731f
C973 avss.t9 dvss 1.2815f
C974 avss.t21 dvss 0.998731f
C975 avss.n222 dvss 0.998731f
C976 avss.n227 dvss 0.177516f
C977 avss.n228 dvss 1.17226f
C978 avss.n229 dvss 0.653412f
C979 avss.n230 dvss 1.44642f
C980 avss.n231 dvss 0.177516f
C981 avss.t25 dvss 0.998731f
C982 avss.t17 dvss 0.998731f
C983 avss.n246 dvss 0.177516f
C984 avss.n247 dvss 0.378264f
C985 avss.n248 dvss 0.401364f
C986 avss.n249 dvss 0.177516f
C987 avss.t80 dvss 0.998731f
C988 avss.t74 dvss 0.998731f
C989 avss.n264 dvss 0.177516f
C990 avss.n265 dvss 1.56554f
C991 avss.n266 dvss 1.24711f
C992 avss.n267 dvss 0.600227f
C993 avss.n268 dvss 1.3851f
C994 avss.t162 dvss 1.73472f
C995 avss.t3 dvss 1.51417f
C996 avss.t136 dvss 1.51417f
C997 avss.t155 dvss 1.51417f
C998 avss.t158 dvss 1.51417f
C999 avss.t141 dvss 1.51417f
C1000 avss.t20 dvss 1.51417f
C1001 avss.t27 dvss 1.5062f
C1002 avss.t95 dvss 1.35433f
C1003 avss.t154 dvss 1.35942f
C1004 avss.t103 dvss 1.35942f
C1005 avss.t85 dvss 1.35942f
C1006 avss.t134 dvss 1.35942f
C1007 avss.t0 dvss 1.35942f
C1008 avss.t66 dvss 1.35942f
C1009 avss.t78 dvss 1.35942f
C1010 avss.t4 dvss 1.35942f
C1011 avss.t119 dvss 1.35942f
C1012 avss.t37 dvss 1.35942f
C1013 avss.t166 dvss 1.36531f
C1014 avss.n269 dvss 1.78687f
C1015 avss.n270 dvss 1.09548f
C1016 avss.n271 dvss 1.35442f
C1017 avss.n272 dvss 14.0235f
C1018 avss.n273 dvss 1.98065f
C1019 avss.t139 dvss 3.05392f
C1020 avss.n274 dvss 1.61326f
C1021 avss.t117 dvss 2.21401f
C1022 avss.n275 dvss 1.96769f
C1023 avss.t43 dvss 1.63078f
C1024 avss.n276 dvss 1.96753f
C1025 avss.t57 dvss 1.63078f
C1026 avss.t61 dvss 1.92756f
C1027 avss.n277 dvss 2.02097f
C1028 avss.n278 dvss 1.57981f
C1029 avss.n279 dvss 0.352908f
C1030 avss.n280 dvss 8.37441f
C1031 avss.n281 dvss 15.798401f
C1032 avss.n282 dvss 2.44293f
C1033 avss.n283 dvss 0.177516f
C1034 avss.n287 dvss 0.289698f
C1035 avss.n289 dvss 0.998731f
C1036 avss.t148 dvss 1.78087f
C1037 avss.t111 dvss 1.99746f
C1038 avss.t58 dvss 1.99746f
C1039 avss.t161 dvss 1.99746f
C1040 avss.t16 dvss 1.48005f
C1041 avss.n291 dvss 0.998731f
C1042 avss.t81 dvss 1.2815f
C1043 avss.t23 dvss 0.998731f
C1044 avss.n294 dvss 0.100238f
C1045 avss.n295 dvss 0.144816f
C1046 avss.n296 dvss 0.136605f
C1047 avss.n298 dvss 0.998731f
C1048 avss.t133 dvss 1.94933f
C1049 avss.t86 dvss 1.27549f
C1050 avss.n299 dvss 1.66809f
C1051 avss.n300 dvss 1.5247f
C1052 avss.n302 dvss 0.158047f
C1053 avss.n303 dvss 0.107219f
C1054 avss.n306 dvss 0.136751f
C1055 avss.t120 dvss 0.569618f
C1056 avss.n312 dvss 0.145184f
C1057 avss.n315 dvss 0.255332f
C1058 avss.n317 dvss 2.87294f
C1059 avss.n318 dvss 0.103631f
C1060 avss.n319 dvss 0.994522f
C1061 avss.n320 dvss 2.53666f
C1062 avss.n321 dvss 5.50604f
C1063 avss.n322 dvss 1.85593f
C1064 avss.t122 dvss 1.4755f
C1065 avss.t38 dvss 1.46417f
C1066 avss.t160 dvss 1.46417f
C1067 avss.t55 dvss 1.46417f
C1068 avss.t32 dvss 0.921721f
C1069 avss.n323 dvss 3.75944f
C1070 avss.n324 dvss 3.81551f
C1071 avss.t100 dvss 0.860352f
C1072 avss.t63 dvss 1.20931f
C1073 avss.t92 dvss 1.07093f
C1074 avss.n325 dvss 0.854336f
C1075 avss.t5 dvss 0.998731f
C1076 avss.n337 dvss 0.177516f
C1077 avss.n338 dvss 1.56743f
C1078 avss.n339 dvss 1.11503f
C1079 avss.n340 dvss 1.80488f
C1080 avss.n341 dvss 6.4046f
C1081 avss.n342 dvss 0.221256f
C1082 avss.n343 dvss 0.134983f
C1083 avss.n344 dvss 0.117108f
C1084 avss.n345 dvss 0.163903f
C1085 avss.n347 dvss 0.998731f
C1086 avss.t45 dvss 1.50411f
C1087 avss.t88 dvss 1.99746f
C1088 avss.t130 dvss 1.99746f
C1089 avss.t118 dvss 2.0755f
C1090 avss.n348 dvss 2.4925f
C1091 avss.n349 dvss 1.1104f
C1092 avss.n350 dvss 0.79897f
C1093 avss.n351 dvss 1.76812f
.ends

