magic
tech sky130A
magscale 1 2
timestamp 1747747376
<< dnwell >>
rect 92 6766 12128 10642
rect 92 3954 9974 6766
rect 92 78 12148 3954
<< nwell >>
rect -24 10436 12244 10758
rect -24 284 298 10436
rect 11922 6972 12244 10436
rect 7118 6034 7988 6713
rect 9768 6650 12244 6972
rect 7118 5356 7372 6034
rect 9768 4070 10090 6650
rect 11613 5041 11667 5393
rect 9768 3748 12264 4070
rect 11942 284 12264 3748
rect -24 -38 12264 284
<< mvnsubdiff >>
rect 49 10665 12171 10685
rect 49 10631 129 10665
rect 12091 10631 12171 10665
rect 49 10611 12171 10631
rect 49 10605 123 10611
rect 49 115 69 10605
rect 103 115 123 10605
rect 12097 10605 12171 10611
rect 12097 6817 12117 10605
rect 12151 6817 12171 10605
rect 12097 6797 12171 6817
rect 9943 6777 12171 6797
rect 9943 6743 10048 6777
rect 12081 6743 12171 6777
rect 9943 6723 12171 6743
rect 9943 6695 10017 6723
rect 9943 4029 9963 6695
rect 9997 4029 10017 6695
rect 9943 3997 10017 4029
rect 9943 3977 12191 3997
rect 9943 3943 10048 3977
rect 12100 3943 12191 3977
rect 9943 3923 12191 3943
rect 49 109 123 115
rect 12117 3909 12191 3923
rect 12117 115 12137 3909
rect 12171 115 12191 3909
rect 12117 109 12191 115
rect 49 89 12191 109
rect 49 55 129 89
rect 12111 55 12191 89
rect 49 35 12191 55
<< mvnsubdiffcont >>
rect 129 10631 12091 10665
rect 69 115 103 10605
rect 12117 6817 12151 10605
rect 10048 6743 12081 6777
rect 9963 4029 9997 6695
rect 10048 3943 12100 3977
rect 12137 115 12171 3909
rect 129 55 12111 89
<< locali >>
rect 62 10665 12153 10670
rect 62 10631 129 10665
rect 12091 10631 12153 10665
rect 62 10605 12153 10631
rect 62 115 69 10605
rect 103 10527 12117 10605
rect 103 7703 186 10527
rect 169 4005 186 7703
rect 295 10315 11944 10429
rect 295 7110 409 10315
rect 11830 7110 11944 10315
rect 295 7091 11944 7110
rect 295 7006 8302 7091
rect 9743 7006 11944 7091
rect 295 6996 11944 7006
rect 12048 9706 12117 10527
rect 12151 10527 12153 10605
rect 12048 7732 12056 9706
rect 496 5313 1636 6996
rect 12048 6893 12117 7732
rect 2181 6751 7885 6752
rect 2134 6725 7885 6751
rect 2134 6668 2219 6725
rect 7862 6668 7885 6725
rect 2134 6593 7885 6668
rect 2134 6150 2288 6593
rect 7565 6151 7885 6593
rect 9855 6866 12117 6893
rect 9855 6841 10031 6866
rect 2134 5924 2503 6150
rect 2777 5924 3119 6150
rect 3393 5924 3735 6150
rect 4009 5924 4351 6150
rect 4625 5924 4967 6150
rect 5241 5924 5583 6150
rect 5857 5924 6199 6150
rect 6473 5924 6815 6150
rect 7565 6150 8009 6151
rect 7089 5924 8009 6150
rect 2134 5469 2288 5924
rect 7881 5469 8009 5924
rect 2134 5312 8009 5469
rect 2181 5311 8009 5312
rect 2181 5310 7900 5311
rect 7877 5206 8000 5207
rect 1020 5047 8000 5206
rect 1020 4611 1151 5047
rect 6591 4618 7453 5047
rect 1020 4449 1122 4611
rect 6591 4607 6796 4618
rect 1278 4605 6796 4607
rect 1278 4448 1661 4605
rect 1916 4448 2217 4605
rect 2472 4448 2773 4605
rect 3028 4448 3329 4605
rect 3584 4448 3885 4605
rect 4140 4448 4441 4605
rect 4696 4448 4997 4605
rect 5252 4448 5553 4605
rect 5808 4448 6109 4605
rect 6364 4449 6796 4605
rect 6952 4607 7453 4618
rect 7877 4607 8000 5047
rect 6952 4449 8000 4607
rect 6364 4448 8000 4449
rect 7877 4013 8000 4448
rect 103 161 186 4005
rect 1131 3963 8000 4013
rect 1131 3928 7905 3963
rect 1131 3873 1183 3928
rect 7858 3873 7905 3928
rect 9855 3943 9880 6841
rect 9945 6801 10031 6841
rect 11457 6817 12117 6866
rect 11457 6801 12151 6817
rect 9945 6777 12151 6801
rect 9945 6743 10048 6777
rect 12081 6743 12151 6777
rect 9945 6731 12151 6743
rect 9945 6695 10004 6731
rect 9945 4029 9963 6695
rect 9997 4029 10004 6695
rect 10519 6573 10924 6580
rect 10519 6444 10633 6573
rect 10519 5942 10924 6444
rect 11596 6250 12049 6252
rect 10193 5734 10924 5942
rect 11591 6249 12049 6250
rect 11591 6122 11623 6249
rect 11827 6122 12049 6249
rect 11591 6119 12049 6122
rect 11591 6023 11734 6119
rect 11591 5960 11616 6023
rect 11723 5960 11734 6023
rect 11591 5797 11734 5960
rect 11591 5767 12049 5797
rect 10452 5491 10924 5734
rect 11593 5722 12049 5767
rect 11593 5540 12049 5615
rect 10188 5476 10924 5491
rect 10188 5475 10813 5476
rect 10188 5248 10231 5475
rect 10404 5248 10813 5475
rect 11595 5396 11738 5540
rect 10188 5234 10813 5248
rect 11572 5388 11738 5396
rect 11572 5192 11601 5388
rect 11735 5192 11738 5388
rect 11572 5131 11738 5192
rect 11572 5057 12054 5131
rect 11576 5056 12054 5057
rect 11257 4826 11577 4957
rect 11624 4939 12054 5014
rect 10217 4685 10423 4687
rect 10217 4683 11590 4685
rect 11624 4683 11739 4939
rect 10217 4673 11739 4683
rect 10217 4513 10231 4673
rect 10408 4637 11739 4673
rect 10408 4513 12054 4637
rect 10217 4498 12054 4513
rect 9945 4017 10004 4029
rect 9945 3977 12171 4017
rect 9945 3943 10048 3977
rect 12100 3943 12171 3977
rect 9855 3909 12171 3943
rect 9855 3893 12137 3909
rect 1131 3854 7905 3873
rect 306 3753 11951 3771
rect 306 3750 5374 3753
rect 306 3671 1862 3750
rect 3521 3674 5374 3750
rect 7033 3674 11951 3753
rect 3521 3671 11951 3674
rect 306 3657 11951 3671
rect 306 3027 420 3657
rect 306 1066 319 3027
rect 413 1066 420 3027
rect 306 409 420 1066
rect 11837 3028 11951 3657
rect 11837 1067 11840 3028
rect 11934 1067 11951 3028
rect 11837 409 11951 1067
rect 306 295 11951 409
rect 12068 161 12137 3893
rect 103 115 12137 161
rect 62 89 12171 115
rect 62 55 129 89
rect 12111 55 12171 89
<< viali >>
rect 88 4005 103 7703
rect 103 4005 169 7703
rect 8302 7006 9743 7091
rect 12056 7732 12117 9706
rect 12117 7732 12144 9706
rect 2219 6668 7862 6725
rect 8319 6547 9723 6880
rect 2503 5924 2777 6151
rect 3119 5924 3393 6151
rect 3735 5924 4009 6151
rect 4351 5924 4625 6151
rect 4967 5924 5241 6151
rect 5583 5924 5857 6151
rect 6199 5924 6473 6151
rect 6815 5924 7089 6151
rect 1122 4442 1278 4611
rect 1661 4448 1916 4605
rect 2217 4448 2472 4605
rect 2773 4448 3028 4605
rect 3329 4448 3584 4605
rect 3885 4448 4140 4605
rect 4441 4448 4696 4605
rect 4997 4448 5252 4605
rect 5553 4448 5808 4605
rect 6109 4448 6364 4605
rect 6796 4449 6952 4618
rect 1183 3873 7858 3928
rect 8312 3923 9716 4256
rect 9880 3943 9945 6841
rect 10031 6801 11457 6866
rect 10633 6444 10929 6573
rect 11623 6122 11827 6249
rect 11616 5960 11723 6023
rect 10231 5248 10404 5475
rect 11601 5192 11735 5388
rect 10231 4513 10408 4673
rect 1862 3671 3521 3750
rect 5374 3674 7033 3753
rect 319 1066 413 3027
rect 11840 1067 11934 3028
<< metal1 >>
rect 514 9788 750 10220
rect 846 9788 1082 10220
rect 1178 9788 1414 10220
rect 1510 9788 1746 10220
rect 1842 9788 2078 10220
rect 2174 9788 2410 10220
rect 2506 9788 2742 10220
rect 2838 9788 3074 10220
rect 3170 9788 3406 10220
rect 3502 9788 3738 10220
rect 3834 9788 4070 10220
rect 4166 9788 4402 10220
rect 4498 9788 4734 10220
rect 4830 9788 5066 10220
rect 5162 9788 5398 10220
rect 5494 9788 5730 10220
rect 5826 9788 6062 10220
rect 6158 9788 6394 10220
rect 6490 9788 6726 10220
rect 6822 9788 7058 10220
rect 7154 9788 7390 10220
rect 7486 9788 7722 10220
rect 7818 9788 8054 10220
rect 8150 9788 8386 10220
rect 8482 9788 8718 10220
rect 8814 9788 9050 10220
rect 9146 9788 9382 10220
rect 9478 9788 9714 10220
rect 9810 9788 10046 10220
rect 10142 9788 10378 10220
rect 10474 9788 10710 10220
rect 10806 9788 11042 10220
rect 11138 9788 11374 10220
rect 11470 9788 11706 10220
rect 12050 9706 12150 9718
rect 12046 7732 12056 9706
rect 12144 7732 12154 9706
rect 12050 7720 12150 7732
rect 82 7703 175 7715
rect 78 4005 88 7703
rect 169 6463 179 7703
rect 513 6641 588 7621
rect 680 7188 916 7620
rect 1012 7188 1248 7620
rect 1344 7188 1580 7620
rect 1676 7188 1912 7620
rect 2008 7188 2244 7620
rect 2340 7188 2576 7620
rect 2672 7188 2908 7620
rect 3004 7188 3240 7620
rect 3336 7188 3572 7620
rect 3668 7188 3904 7620
rect 4000 7188 4236 7620
rect 4332 7188 4568 7620
rect 4664 7188 4900 7620
rect 4996 7188 5232 7620
rect 5328 7188 5564 7620
rect 5660 7188 5896 7620
rect 5992 7188 6228 7620
rect 6324 7188 6560 7620
rect 6656 7188 6892 7620
rect 6988 7188 7224 7620
rect 7320 7188 7556 7620
rect 7652 7188 7888 7620
rect 7984 7188 8220 7620
rect 8316 7188 8552 7620
rect 8648 7188 8884 7620
rect 8980 7188 9216 7620
rect 9312 7188 9548 7620
rect 9644 7188 9880 7620
rect 9976 7188 10212 7620
rect 10308 7188 10544 7620
rect 10640 7188 10876 7620
rect 10972 7188 11208 7620
rect 11304 7188 11540 7620
rect 627 7100 1828 7103
rect 8285 7100 9768 7110
rect 627 7091 9768 7100
rect 627 7089 8302 7091
rect 627 6962 654 7089
rect 1795 7006 8302 7089
rect 9743 7006 9768 7091
rect 1795 6962 9768 7006
rect 627 6945 9768 6962
rect 807 6944 9768 6945
rect 8172 6924 9768 6944
rect 8285 6901 9768 6924
rect 9837 7019 11494 7044
rect 9837 6901 9877 7019
rect 11458 6901 11494 7019
rect 8285 6880 9767 6901
rect 2137 6818 7913 6848
rect 2137 6753 2190 6818
rect 7886 6753 7913 6818
rect 2137 6725 7913 6753
rect 2137 6668 2219 6725
rect 7862 6668 7913 6725
rect 2137 6658 7913 6668
rect 513 6590 1839 6641
rect 169 5310 1632 6463
rect 169 4005 179 5310
rect 1439 4946 1449 4967
rect 1194 4623 1278 4871
rect 1348 4720 1376 4937
rect 1384 4906 1449 4946
rect 1439 4905 1449 4906
rect 1606 4905 1616 4967
rect 1116 4611 1284 4623
rect 1112 4442 1122 4611
rect 1278 4442 1288 4611
rect 1116 4430 1284 4442
rect 1454 4129 1486 4868
rect 1788 4790 1839 6590
rect 8285 6547 8319 6880
rect 9723 6547 9767 6880
rect 2373 6475 6862 6522
rect 8285 6506 9767 6547
rect 9837 6866 11494 6901
rect 9837 6841 10031 6866
rect 2373 5696 2420 6475
rect 2483 6265 2514 6475
rect 2573 6157 2673 6415
rect 2491 6151 2789 6157
rect 2491 5924 2503 6151
rect 2777 5924 2789 6151
rect 2491 5918 2789 5924
rect 2336 5649 2420 5696
rect 1960 5063 1970 5084
rect 1903 5022 1970 5063
rect 2127 5063 2137 5084
rect 2127 5026 2217 5063
rect 2127 5022 2137 5026
rect 1903 4722 1940 5022
rect 1649 4605 1928 4611
rect 1649 4448 1661 4605
rect 1916 4448 1928 4605
rect 1649 4442 1928 4448
rect 1747 4185 1831 4442
rect 1904 4129 1937 4328
rect 2009 4129 2049 4879
rect 2180 4752 2217 5026
rect 2336 4786 2383 5649
rect 2482 5088 2514 5802
rect 2588 5652 2692 5918
rect 2985 5653 3029 6422
rect 3099 6265 3130 6475
rect 3189 6157 3289 6415
rect 3107 6151 3405 6157
rect 3107 5924 3119 6151
rect 3393 5924 3405 6151
rect 3107 5918 3405 5924
rect 3092 5328 3131 5807
rect 2993 5163 3003 5328
rect 3060 5286 3131 5328
rect 3190 5516 3229 5734
rect 3601 5653 3645 6422
rect 3715 6265 3746 6475
rect 3805 6157 3905 6415
rect 3723 6151 4021 6157
rect 3723 5924 3735 6151
rect 4009 5924 4021 6151
rect 3723 5918 4021 5924
rect 3190 5426 3204 5516
rect 3414 5426 3424 5516
rect 3190 5326 3229 5426
rect 3708 5326 3747 5807
rect 3190 5287 3747 5326
rect 3819 5516 3858 5738
rect 4217 5653 4261 6422
rect 4331 6265 4362 6475
rect 4421 6157 4521 6415
rect 4339 6151 4637 6157
rect 4339 5924 4351 6151
rect 4625 5924 4637 6151
rect 4339 5918 4637 5924
rect 3819 5426 3835 5516
rect 4045 5426 4055 5516
rect 3819 5328 3858 5426
rect 4324 5328 4363 5807
rect 3819 5289 4363 5328
rect 4445 5516 4484 5745
rect 4833 5653 4877 6422
rect 4947 6265 4978 6475
rect 5037 6157 5137 6415
rect 4955 6151 5253 6157
rect 4955 5924 4967 6151
rect 5241 5924 5253 6151
rect 4955 5918 5253 5924
rect 4445 5426 4467 5516
rect 4677 5426 4687 5516
rect 4445 5328 4484 5426
rect 4940 5328 4979 5807
rect 4445 5289 4979 5328
rect 5048 5516 5087 5737
rect 5449 5653 5493 6422
rect 5563 6265 5594 6475
rect 5653 6157 5753 6415
rect 5571 6151 5869 6157
rect 5571 5924 5583 6151
rect 5857 5924 5869 6151
rect 5571 5918 5869 5924
rect 5048 5426 5071 5516
rect 5281 5426 5291 5516
rect 5048 5328 5087 5426
rect 5556 5328 5595 5807
rect 5048 5289 5595 5328
rect 5672 5498 5711 5744
rect 6065 5653 6109 6422
rect 6179 6265 6210 6475
rect 6269 6157 6369 6415
rect 6187 6151 6485 6157
rect 6187 5924 6199 6151
rect 6473 5924 6485 6151
rect 6187 5918 6485 5924
rect 5874 5498 5884 5516
rect 5672 5442 5884 5498
rect 5672 5328 5711 5442
rect 5874 5426 5884 5442
rect 6094 5426 6104 5516
rect 6172 5328 6211 5807
rect 5672 5289 6211 5328
rect 6283 5328 6322 5741
rect 6681 5653 6725 6422
rect 6795 6265 6826 6475
rect 6885 6157 6985 6415
rect 7502 6173 7512 6272
rect 7872 6173 7882 6272
rect 6803 6151 7101 6157
rect 6803 5924 6815 6151
rect 7089 5924 7101 6151
rect 6803 5918 7101 5924
rect 6788 5328 6827 5807
rect 6905 5332 6944 5744
rect 7511 5666 7595 6173
rect 8020 5967 8030 5988
rect 7758 5929 8030 5967
rect 7656 5513 7700 5824
rect 7203 5469 7700 5513
rect 6283 5289 6827 5328
rect 3060 5163 3070 5286
rect 2472 5026 2482 5088
rect 2639 5026 2649 5088
rect 2459 4752 2496 4959
rect 2180 4715 2496 4752
rect 2205 4605 2484 4611
rect 2205 4448 2217 4605
rect 2472 4448 2484 4605
rect 2205 4442 2484 4448
rect 2303 4431 2395 4442
rect 2311 4188 2395 4431
rect 2461 4130 2494 4333
rect 2561 4188 2603 4877
rect 2904 4681 2946 4874
rect 3016 4720 3055 5163
rect 3190 5015 3229 5287
rect 3128 4976 3229 5015
rect 3128 4787 3167 4976
rect 3460 4681 3502 4874
rect 3572 4720 3611 5287
rect 3819 5016 3858 5289
rect 3679 4977 3858 5016
rect 3679 4781 3718 4977
rect 4016 4681 4058 4874
rect 4128 4720 4167 5289
rect 4445 5018 4484 5289
rect 4235 4979 4484 5018
rect 4235 4789 4274 4979
rect 4572 4681 4614 4874
rect 4684 4720 4723 5289
rect 5048 5021 5087 5289
rect 4789 4982 5087 5021
rect 4789 4781 4828 4982
rect 5128 4681 5170 4874
rect 5240 4720 5279 5289
rect 5672 5020 5711 5289
rect 5347 4981 5711 5020
rect 5347 4782 5386 4981
rect 5684 4681 5726 4874
rect 5796 4720 5835 5289
rect 6283 5027 6322 5289
rect 5910 4988 6322 5027
rect 5910 4786 5949 4988
rect 6240 4681 6282 4874
rect 6352 4720 6391 5289
rect 6892 5167 6902 5332
rect 6959 5290 6969 5332
rect 7203 5290 7247 5469
rect 6959 5223 7247 5290
rect 6959 5167 6969 5223
rect 6905 5032 6944 5167
rect 6457 4993 6944 5032
rect 6457 4787 6496 4993
rect 2904 4639 3159 4681
rect 3460 4639 3715 4681
rect 4016 4639 4271 4681
rect 4572 4639 4827 4681
rect 5128 4639 5383 4681
rect 5684 4639 5939 4681
rect 6240 4639 6495 4681
rect 2761 4605 3040 4611
rect 2761 4448 2773 4605
rect 3028 4448 3040 4605
rect 2761 4442 3040 4448
rect 2859 4431 2951 4442
rect 2867 4188 2951 4431
rect 3017 4130 3050 4333
rect 3117 4188 3159 4639
rect 3317 4605 3596 4611
rect 3317 4448 3329 4605
rect 3584 4448 3596 4605
rect 3317 4442 3596 4448
rect 3415 4431 3507 4442
rect 3423 4188 3507 4431
rect 3573 4130 3606 4333
rect 3673 4188 3715 4639
rect 3873 4605 4152 4611
rect 3873 4448 3885 4605
rect 4140 4448 4152 4605
rect 3873 4442 4152 4448
rect 3971 4431 4063 4442
rect 3979 4188 4063 4431
rect 4129 4130 4162 4333
rect 4229 4188 4271 4639
rect 4429 4605 4708 4611
rect 4429 4448 4441 4605
rect 4696 4448 4708 4605
rect 4429 4442 4708 4448
rect 4527 4431 4619 4442
rect 4535 4188 4619 4431
rect 4685 4130 4718 4333
rect 4785 4188 4827 4639
rect 4985 4605 5264 4611
rect 4985 4448 4997 4605
rect 5252 4448 5264 4605
rect 4985 4442 5264 4448
rect 5083 4431 5175 4442
rect 5091 4188 5175 4431
rect 5241 4130 5274 4333
rect 5341 4188 5383 4639
rect 5541 4605 5820 4611
rect 5541 4448 5553 4605
rect 5808 4448 5820 4605
rect 5541 4442 5820 4448
rect 5639 4431 5731 4442
rect 5647 4188 5731 4431
rect 5797 4130 5830 4333
rect 5897 4188 5939 4639
rect 6097 4605 6376 4611
rect 6097 4448 6109 4605
rect 6364 4448 6376 4605
rect 6097 4442 6376 4448
rect 6195 4431 6287 4442
rect 6203 4188 6287 4431
rect 6353 4130 6386 4333
rect 6453 4188 6495 4639
rect 6790 4618 6958 4630
rect 6790 4613 6796 4618
rect 6656 4605 6796 4613
rect 6656 4448 6665 4605
rect 6952 4449 6958 4618
rect 6920 4448 6958 4449
rect 6656 4439 6958 4448
rect 6790 4437 6958 4439
rect 7203 4447 7247 5223
rect 7544 4623 7582 4860
rect 7649 4743 7685 4933
rect 7758 4785 7796 5929
rect 8020 5910 8030 5929
rect 8221 5910 8231 5988
rect 8050 5145 8329 5179
rect 8050 4961 8084 5145
rect 7930 4897 7940 4961
rect 8127 4897 8137 4961
rect 7649 4707 8069 4743
rect 8033 4638 8069 4707
rect 7544 4585 7795 4623
rect 8033 4599 8097 4638
rect 6824 4274 6908 4437
rect 7203 4404 7690 4447
rect 7261 4403 7690 4404
rect 6824 4273 7584 4274
rect 6824 4191 7594 4273
rect 6824 4190 7482 4191
rect 1454 4081 6404 4129
rect 7646 4124 7690 4403
rect 7757 4190 7795 4585
rect 8087 4574 8097 4599
rect 8284 4574 8294 4638
rect 9837 4316 9880 6841
rect 9725 4306 9880 4316
rect 8268 4256 9880 4306
rect 82 3993 175 4005
rect 1129 3928 7903 4013
rect 1129 3873 1183 3928
rect 7858 3873 7903 3928
rect 8268 3923 8312 4256
rect 9716 3943 9880 4256
rect 9945 6801 10031 6841
rect 11457 6801 11494 6866
rect 9945 6774 11494 6801
rect 9945 3943 10014 6774
rect 11658 6702 11733 7627
rect 10494 6627 11733 6702
rect 10267 6483 10277 6555
rect 10453 6483 10463 6555
rect 10254 5988 10307 6188
rect 10391 6102 10453 6483
rect 10065 5916 10075 5988
rect 10251 5934 10307 5988
rect 10251 5916 10261 5934
rect 10352 5780 10384 6064
rect 10240 5708 10250 5780
rect 10426 5708 10436 5780
rect 10352 5641 10384 5643
rect 10212 5569 10222 5641
rect 10398 5569 10408 5641
rect 10217 5475 10423 5493
rect 10217 5248 10231 5475
rect 10404 5248 10423 5475
rect 10217 4673 10423 5248
rect 10217 4513 10231 4673
rect 10408 4513 10423 4673
rect 10217 4500 10423 4513
rect 10494 4131 10569 6627
rect 10621 6573 10941 6579
rect 10621 6444 10633 6573
rect 10929 6444 10941 6573
rect 11864 6564 12244 7141
rect 10621 6438 10941 6444
rect 11142 6554 12244 6564
rect 11142 6455 11153 6554
rect 11513 6455 12244 6554
rect 11142 6364 12244 6455
rect 10638 6177 10648 6276
rect 11008 6177 11018 6276
rect 11142 6249 11839 6364
rect 10644 4934 10806 6177
rect 11142 6122 11623 6249
rect 11827 6122 11839 6249
rect 11142 6116 11839 6122
rect 11142 6039 11629 6116
rect 11142 6023 11838 6039
rect 11142 5960 11616 6023
rect 11723 5960 11838 6023
rect 11142 5945 11838 5960
rect 11142 5943 11342 5945
rect 11829 5944 11838 5945
rect 11938 5938 11986 6044
rect 11938 5890 12060 5938
rect 11818 5829 11904 5883
rect 11489 5655 11499 5672
rect 11428 5600 11499 5655
rect 11675 5663 11685 5672
rect 11818 5663 11859 5829
rect 11675 5614 11859 5663
rect 11675 5600 11685 5614
rect 11428 5290 11466 5600
rect 11818 5431 11859 5614
rect 11887 5613 11897 5782
rect 11966 5613 11976 5782
rect 11910 5530 11976 5613
rect 11595 5388 11741 5400
rect 11338 5252 11466 5290
rect 11338 5136 11376 5252
rect 11503 5222 11601 5388
rect 11435 5192 11601 5222
rect 11735 5192 11841 5388
rect 11435 5190 11841 5192
rect 11435 5180 11741 5190
rect 11435 5140 11715 5180
rect 11253 5026 11263 5098
rect 11439 5026 11449 5098
rect 11503 4934 11715 5140
rect 11935 5127 11976 5530
rect 10644 4734 11715 4934
rect 11787 5086 11976 5127
rect 11787 4786 11828 5086
rect 12012 5038 12060 5890
rect 11939 4990 12060 5038
rect 11939 4786 11987 4990
rect 11155 4391 11715 4734
rect 11777 4671 11787 4730
rect 11973 4671 11983 4730
rect 11155 4191 12264 4391
rect 10494 4056 11733 4131
rect 9716 3923 10014 3943
rect 8268 3892 10014 3923
rect 1129 3856 7903 3873
rect 1850 3750 3533 3756
rect 1850 3671 1862 3750
rect 3521 3671 3533 3750
rect 1850 3665 3533 3671
rect 5362 3753 7045 3759
rect 5362 3674 5374 3753
rect 7033 3674 7045 3753
rect 5362 3668 7045 3674
rect 62 3525 4256 3532
rect 62 3116 76 3525
rect 351 3116 4256 3525
rect 62 3100 4256 3116
rect 4352 3100 4588 3532
rect 4684 3100 4920 3532
rect 5016 3100 5252 3532
rect 5348 3100 5584 3532
rect 5680 3100 5916 3532
rect 6012 3100 6248 3532
rect 6344 3100 6580 3532
rect 6676 3100 6912 3532
rect 7008 3100 7244 3532
rect 7340 3100 7576 3532
rect 7672 3100 7908 3532
rect 8004 3100 8240 3532
rect 8336 3100 8572 3532
rect 8668 3100 8904 3532
rect 9000 3100 9236 3532
rect 9332 3100 9568 3532
rect 9664 3100 9900 3532
rect 9996 3100 10232 3532
rect 10328 3100 10564 3532
rect 10660 3100 10896 3532
rect 10992 3100 11228 3532
rect 11324 3100 11560 3532
rect 313 3027 419 3039
rect 309 1066 319 3027
rect 413 1066 423 3027
rect 313 1054 419 1066
rect 522 932 716 3100
rect 11658 3097 11733 4056
rect 11864 3616 12264 4191
rect 11834 3028 11940 3040
rect 11830 1067 11840 3028
rect 11934 1067 11944 3028
rect 11834 1055 11940 1067
rect 522 930 770 932
rect 866 930 1102 932
rect 1198 930 1434 932
rect 1530 930 1766 932
rect 1862 930 2098 932
rect 2194 930 2430 932
rect 2526 930 2762 932
rect 2858 930 3094 932
rect 3190 930 3426 932
rect 3522 930 3758 932
rect 3854 930 4090 932
rect 522 498 4092 930
rect 4186 500 4422 932
rect 4518 500 4754 932
rect 4850 500 5086 932
rect 5182 500 5418 932
rect 5514 500 5750 932
rect 5846 500 6082 932
rect 6178 500 6414 932
rect 6510 500 6746 932
rect 6842 500 7078 932
rect 7174 500 7410 932
rect 7506 500 7742 932
rect 7838 500 8074 932
rect 8170 500 8406 932
rect 8502 500 8738 932
rect 8834 500 9070 932
rect 9166 500 9402 932
rect 9498 500 9734 932
rect 9830 500 10066 932
rect 10162 500 10398 932
rect 10494 500 10730 932
rect 10826 500 11062 932
rect 11158 500 11394 932
rect 11490 500 11726 932
<< via1 >>
rect 12056 7732 12144 9706
rect 88 4005 169 7703
rect 654 6962 1795 7089
rect 9877 6901 11458 7019
rect 2190 6753 7886 6818
rect 1449 4905 1606 4967
rect 1122 4442 1278 4611
rect 8319 6547 9723 6880
rect 2503 5924 2777 6151
rect 1970 5022 2127 5084
rect 1661 4448 1916 4605
rect 3119 5924 3393 6151
rect 3003 5163 3060 5328
rect 3735 5924 4009 6151
rect 3204 5426 3414 5516
rect 4351 5924 4625 6151
rect 3835 5426 4045 5516
rect 4967 5924 5241 6151
rect 4467 5426 4677 5516
rect 5583 5924 5857 6151
rect 5071 5426 5281 5516
rect 6199 5924 6473 6151
rect 5884 5426 6094 5516
rect 7512 6173 7872 6272
rect 6815 5924 7089 6151
rect 2482 5026 2639 5088
rect 2217 4448 2472 4605
rect 6902 5167 6959 5332
rect 2773 4448 3028 4605
rect 3329 4448 3584 4605
rect 3885 4448 4140 4605
rect 4441 4448 4696 4605
rect 4997 4448 5252 4605
rect 5553 4448 5808 4605
rect 6109 4448 6364 4605
rect 6665 4449 6796 4605
rect 6796 4449 6920 4605
rect 6665 4448 6920 4449
rect 8030 5910 8221 5988
rect 7940 4897 8127 4961
rect 8097 4574 8284 4638
rect 1183 3873 7858 3928
rect 8312 3923 9716 4256
rect 10277 6483 10453 6555
rect 10075 5916 10251 5988
rect 10250 5708 10426 5780
rect 10222 5569 10398 5641
rect 10633 6444 10929 6573
rect 11153 6455 11513 6554
rect 10648 6177 11008 6276
rect 11499 5600 11675 5672
rect 11897 5613 11966 5782
rect 11263 5026 11439 5098
rect 11787 4671 11973 4730
rect 1862 3671 3521 3750
rect 5374 3674 7033 3753
rect 76 3116 351 3525
rect 319 1066 413 3027
rect 11840 1067 11934 3028
<< metal2 >>
rect 12056 9715 12144 9716
rect -24 9706 12244 9715
rect -24 7732 12056 9706
rect 12144 7732 12244 9706
rect -24 7721 12244 7732
rect 68 7703 358 7721
rect 68 4005 88 7703
rect 169 4005 358 7703
rect 627 7089 1828 7103
rect 627 7085 654 7089
rect 68 3525 358 4005
rect 68 3116 76 3525
rect 351 3116 358 3525
rect 68 3110 358 3116
rect 625 6962 654 7085
rect 1795 6962 1828 7089
rect 625 6945 1828 6962
rect 625 6464 1175 6945
rect 2453 6865 4111 7721
rect 5409 6865 7067 7721
rect 8285 6901 9768 7110
rect 9837 7019 11494 7721
rect 9837 6901 9877 7019
rect 11458 6901 11494 7019
rect 8285 6880 9767 6901
rect 9837 6882 11494 6901
rect 2119 6818 7954 6865
rect 2119 6753 2190 6818
rect 7886 6753 7954 6818
rect 2119 6655 7954 6753
rect 625 5307 1635 6464
rect 2453 6199 4111 6655
rect 5409 6199 7067 6655
rect 8285 6547 8319 6880
rect 9723 6547 9767 6880
rect 10633 6574 10929 6583
rect 8285 6506 9767 6547
rect 10263 6573 11518 6574
rect 10263 6555 10633 6573
rect 10263 6483 10277 6555
rect 10453 6483 10633 6555
rect 10263 6444 10633 6483
rect 10929 6554 11518 6573
rect 10929 6455 11153 6554
rect 11513 6455 11518 6554
rect 10929 6444 11518 6455
rect 10263 6442 11518 6444
rect 10633 6434 10929 6442
rect 7512 6274 7872 6282
rect 10648 6276 11008 6286
rect 7512 6272 10648 6274
rect 2131 6151 7166 6199
rect 7872 6177 10648 6272
rect 7872 6176 11008 6177
rect 7512 6163 7872 6173
rect 10648 6167 11008 6176
rect 2131 5924 2503 6151
rect 2777 5924 3119 6151
rect 3393 5924 3735 6151
rect 4009 5924 4351 6151
rect 4625 5924 4967 6151
rect 5241 5924 5583 6151
rect 5857 5924 6199 6151
rect 6473 5924 6815 6151
rect 7089 5924 7166 6151
rect 2131 5883 7166 5924
rect 8030 5988 8221 5998
rect 10075 5988 10251 5998
rect 8221 5929 9972 5973
rect 10074 5929 10075 5973
rect 8030 5900 8221 5910
rect 9928 5876 9972 5929
rect 10251 5929 11574 5973
rect 10075 5906 10251 5916
rect 9928 5832 11424 5876
rect 10250 5780 10426 5790
rect 10250 5698 10426 5708
rect 11380 5654 11424 5832
rect 11530 5759 11574 5929
rect 11897 5782 11966 5792
rect 11530 5715 11897 5759
rect 11499 5672 11675 5682
rect 10222 5641 10398 5651
rect 2521 5592 2619 5602
rect 3587 5592 3685 5602
rect 3204 5523 3414 5526
rect 2619 5516 3414 5523
rect 2619 5457 3204 5516
rect 2521 5426 3204 5457
rect 2521 5418 3414 5426
rect 2521 5367 2619 5418
rect 3204 5416 3414 5418
rect 4653 5592 4751 5602
rect 3685 5526 3851 5527
rect 3685 5516 4045 5526
rect 3685 5457 3835 5516
rect 3587 5426 3835 5457
rect 3587 5417 4045 5426
rect 3587 5367 3685 5417
rect 3835 5416 4045 5417
rect 4467 5516 4653 5526
rect 5719 5592 5817 5602
rect 4677 5426 4751 5457
rect 4467 5416 4751 5426
rect 5071 5516 5719 5526
rect 5281 5457 5719 5516
rect 6785 5592 6883 5602
rect 6082 5526 6785 5527
rect 5281 5426 5817 5457
rect 5071 5417 5817 5426
rect 5071 5416 5281 5417
rect 4653 5367 4751 5416
rect 5719 5367 5817 5417
rect 5884 5516 6785 5526
rect 6094 5457 6785 5516
rect 6094 5426 6883 5457
rect 5884 5417 6883 5426
rect 5884 5416 6094 5417
rect 6785 5367 6883 5417
rect 3003 5328 3060 5338
rect 625 4644 1175 5307
rect 6902 5332 6959 5342
rect 3060 5220 6902 5261
rect 3003 5153 3060 5163
rect 6902 5157 6959 5167
rect 1970 5084 2127 5094
rect 2482 5088 2639 5098
rect 1932 5023 1970 5084
rect 2127 5026 2482 5084
rect 2639 5026 8263 5084
rect 2127 5023 8263 5026
rect 1970 5012 2127 5022
rect 2482 5016 2639 5023
rect 1449 4967 1606 4977
rect 7930 4961 8127 4971
rect 7930 4950 7940 4961
rect 1606 4905 7940 4950
rect 1449 4895 1606 4905
rect 7940 4887 8127 4897
rect 8202 4926 8263 5023
rect 8202 4865 8538 4926
rect 625 4611 7135 4644
rect 8097 4639 8284 4648
rect 9688 4639 9753 5600
rect 11380 5610 11499 5654
rect 12042 5759 12242 5830
rect 11966 5715 12242 5759
rect 12042 5630 12242 5715
rect 11897 5603 11966 5613
rect 11499 5590 11675 5600
rect 10222 5559 10398 5569
rect 11016 5391 11569 5445
rect 11263 5098 11439 5108
rect 11515 5086 11569 5391
rect 11439 5039 11569 5086
rect 11263 5016 11439 5026
rect 11515 4913 11569 5039
rect 12042 4913 12242 4986
rect 11515 4859 12242 4913
rect 11854 4740 11910 4859
rect 12042 4786 12242 4859
rect 11787 4730 11973 4740
rect 11787 4661 11973 4671
rect 625 4442 1122 4611
rect 1278 4605 7135 4611
rect 1278 4448 1661 4605
rect 1916 4448 2217 4605
rect 2472 4448 2773 4605
rect 3028 4448 3329 4605
rect 3584 4448 3885 4605
rect 4140 4448 4441 4605
rect 4696 4448 4997 4605
rect 5252 4448 5553 4605
rect 5808 4448 6109 4605
rect 6364 4448 6665 4605
rect 6920 4448 7135 4605
rect 8095 4638 9753 4639
rect 8095 4574 8097 4638
rect 8284 4574 9753 4638
rect 8097 4564 8284 4574
rect 1278 4442 7135 4448
rect 625 4342 7135 4442
rect 625 4038 1175 4342
rect 1861 4038 3520 4342
rect 5375 4038 7034 4342
rect 8268 4256 9750 4306
rect 625 3928 7930 4038
rect 625 3873 1183 3928
rect 7858 3873 7930 3928
rect 8268 3923 8312 4256
rect 9716 3923 9750 4256
rect 8268 3892 9750 3923
rect 625 3824 7930 3873
rect 625 3044 1175 3824
rect 1861 3750 3521 3824
rect 1861 3671 1862 3750
rect 1861 3661 3521 3671
rect 5374 3753 7034 3824
rect 7033 3674 7034 3753
rect 5374 3664 7034 3674
rect 1861 3044 3520 3661
rect 5375 3044 7034 3664
rect -24 3028 12264 3044
rect -24 3027 11840 3028
rect -24 1066 319 3027
rect 413 2990 11840 3027
rect 413 2723 3091 2990
rect 7477 2723 11840 2990
rect 413 1067 11840 2723
rect 11934 1067 12264 3028
rect 413 1066 12264 1067
rect -24 1050 12264 1066
<< via2 >>
rect 2521 5457 2619 5592
rect 3587 5457 3685 5592
rect 4653 5516 4751 5592
rect 4653 5457 4677 5516
rect 4677 5457 4751 5516
rect 5719 5457 5817 5592
rect 6785 5457 6883 5592
rect 3091 2723 7477 2990
<< metal3 >>
rect 2511 5672 2629 5677
rect 2511 5457 2521 5672
rect 2619 5457 2629 5672
rect 2511 5452 2629 5457
rect 3577 5672 3695 5677
rect 3577 5457 3587 5672
rect 3685 5457 3695 5672
rect 3577 5452 3695 5457
rect 4643 5672 4761 5677
rect 4643 5457 4653 5672
rect 4751 5457 4761 5672
rect 4643 5452 4761 5457
rect 5709 5672 5827 5677
rect 5709 5457 5719 5672
rect 5817 5457 5827 5672
rect 5709 5452 5827 5457
rect 6775 5672 6893 5677
rect 6775 5457 6785 5672
rect 6883 5457 6893 5672
rect 6775 5452 6893 5457
rect 3204 3930 3298 5210
rect 4270 3930 4364 5210
rect 5336 3931 5430 5211
rect 6402 3931 6496 5211
rect 3094 3453 3104 3703
rect 3202 3453 3212 3703
rect 3094 2995 3212 3453
rect 4160 3453 4170 3703
rect 4268 3453 4278 3703
rect 4160 2995 4278 3453
rect 5226 3453 5236 3703
rect 5334 3453 5344 3703
rect 5226 2995 5344 3453
rect 6292 3453 6302 3703
rect 6400 3453 6410 3703
rect 6292 2995 6410 3453
rect 7358 3453 7368 3703
rect 7466 3453 7476 3703
rect 7358 2995 7476 3453
rect 3081 2990 7487 2995
rect 3081 2723 3091 2990
rect 7477 2723 7487 2990
rect 3081 2718 7487 2723
<< via3 >>
rect 2521 5592 2619 5672
rect 2521 5457 2619 5592
rect 3587 5592 3685 5672
rect 3587 5457 3685 5592
rect 4653 5592 4751 5672
rect 4653 5457 4751 5592
rect 5719 5592 5817 5672
rect 5719 5457 5817 5592
rect 6785 5592 6883 5672
rect 6785 5457 6883 5592
rect 3104 3453 3202 3703
rect 4170 3453 4268 3703
rect 5236 3453 5334 3703
rect 6302 3453 6400 3703
rect 7368 3453 7466 3703
<< metal4 >>
rect 2510 5672 2630 5678
rect 2510 5457 2521 5672
rect 2619 5457 2630 5672
rect 2510 5450 2630 5457
rect 3576 5672 3696 5678
rect 3576 5457 3587 5672
rect 3685 5457 3696 5672
rect 3576 5450 3696 5457
rect 4642 5672 4762 5678
rect 4642 5457 4653 5672
rect 4751 5457 4762 5672
rect 4642 5450 4762 5457
rect 5708 5672 5828 5678
rect 5708 5457 5719 5672
rect 5817 5457 5828 5672
rect 5708 5450 5828 5457
rect 6774 5672 6894 5678
rect 6774 5457 6785 5672
rect 6883 5457 6894 5672
rect 6774 5450 6894 5457
rect 2521 4328 2619 5450
rect 3587 4328 3685 5450
rect 4653 4328 4751 5450
rect 5719 4328 5817 5450
rect 6785 4328 6883 5450
rect 3104 3704 3202 4080
rect 4170 3704 4268 4080
rect 5236 3704 5334 4080
rect 6302 3704 6400 4080
rect 7368 3704 7466 4080
rect 3103 3703 3203 3704
rect 3103 3453 3104 3703
rect 3202 3453 3203 3703
rect 3103 3452 3203 3453
rect 4169 3703 4269 3704
rect 4169 3453 4170 3703
rect 4268 3453 4269 3703
rect 4169 3452 4269 3453
rect 5235 3703 5335 3704
rect 5235 3453 5236 3703
rect 5334 3453 5335 3703
rect 5235 3452 5335 3453
rect 6301 3703 6401 3704
rect 6301 3453 6302 3703
rect 6400 3453 6401 3703
rect 6301 3452 6401 3453
rect 7367 3703 7467 3704
rect 7367 3453 7368 3703
rect 7466 3453 7467 3703
rect 7367 3452 7467 3453
use sky130_fd_pr__diode_pw2nd_05v5_FT76RJ  D3 paramcells
timestamp 1747747376
transform 1 0 10339 0 1 5604
box -183 -183 183 183
use rc_osc_level_shifter  rc_osc_level_shifter_0
timestamp 1747747376
transform -1 0 10932 0 -1 4214
box -422 -2544 2736 144
use sky130_fd_pr__cap_mim_m3_1_AZFCP3  sky130_fd_pr__cap_mim_m3_1_AZFCP3_1 paramcells
timestamp 1747747376
transform 1 0 6982 0 1 4571
box -486 -640 486 640
use sky130_fd_pr__nfet_01v8_L9WNCD  sky130_fd_pr__nfet_01v8_L9WNCD_0 paramcells
timestamp 1747747376
transform 1 0 11875 0 1 5958
box -211 -229 211 229
use sky130_fd_pr__pfet_01v8_2Z69BZ  sky130_fd_pr__pfet_01v8_2Z69BZ_0 paramcells
timestamp 1747747376
transform 1 0 11402 0 1 5145
box -211 -226 211 226
use sky130_fd_pr__pfet_01v8_LGS3BL  sky130_fd_pr__pfet_01v8_LGS3BL_0 paramcells
timestamp 1747747376
transform 1 0 11878 0 -1 5325
box -211 -284 211 284
use sky130_fd_pr__res_xhigh_po_0p35_DEAPHQ  sky130_fd_pr__res_xhigh_po_0p35_DEAPHQ_0 paramcells
timestamp 1747747376
transform 1 0 6130 0 1 2016
box -5762 -1682 5762 1682
use sky130_fd_pr__res_xhigh_po_0p35_DEAPHQ  sky130_fd_pr__res_xhigh_po_0p35_DEAPHQ_1
timestamp 1747747376
transform 1 0 6110 0 1 8704
box -5762 -1682 5762 1682
use sky130_fd_pr__cap_mim_m3_1_AZFCP3  XC1
timestamp 1747747376
transform 1 0 2718 0 1 4570
box -486 -640 486 640
use sky130_fd_pr__cap_mim_m3_1_AZFCP3  XC2
timestamp 1747747376
transform 1 0 3784 0 1 4570
box -486 -640 486 640
use sky130_fd_pr__cap_mim_m3_1_AZFCP3  XC3
timestamp 1747747376
transform 1 0 4850 0 1 4571
box -486 -640 486 640
use sky130_fd_pr__cap_mim_m3_1_AZFCP3  XC4
timestamp 1747747376
transform 1 0 5916 0 1 4571
box -486 -640 486 640
use sky130_fd_pr__nfet_g5v0d10v5_6XHUDR  XM1 paramcells
timestamp 1747747376
transform 1 0 3032 0 1 4830
box -278 -300 278 300
use sky130_fd_pr__pfet_g5v0d10v5_6ELFTH  XM2 paramcells
timestamp 1747747376
transform 1 0 3114 0 1 5695
box -308 -339 308 339
use sky130_fd_pr__pfet_g5v0d10v5_6ELFTH  XM3
timestamp 1747747376
transform 1 0 3730 0 1 5695
box -308 -339 308 339
use sky130_fd_pr__nfet_g5v0d10v5_6XHUDR  XM4
timestamp 1747747376
transform 1 0 3588 0 1 4830
box -278 -300 278 300
use sky130_fd_pr__nfet_01v8_L9WNCD  XM5
timestamp 1747747376
transform 1 0 11882 0 1 4794
box -211 -229 211 229
use sky130_fd_pr__pfet_g5v0d10v5_6ELFTH  XM7
timestamp 1747747376
transform 1 0 4962 0 1 5695
box -308 -339 308 339
use sky130_fd_pr__nfet_g5v0d10v5_6XHUDR  XM8
timestamp 1747747376
transform 1 0 4700 0 1 4830
box -278 -300 278 300
use sky130_fd_pr__pfet_g5v0d10v5_6ELFTH  XM9
timestamp 1747747376
transform 1 0 4346 0 1 5695
box -308 -339 308 339
use sky130_fd_pr__nfet_g5v0d10v5_6XHUDR  XM10
timestamp 1747747376
transform 1 0 4144 0 1 4830
box -278 -300 278 300
use sky130_fd_pr__pfet_g5v0d10v5_6ELFTH  XM11
timestamp 1747747376
transform 1 0 7680 0 1 5695
box -308 -339 308 339
use sky130_fd_pr__nfet_g5v0d10v5_6XHUDR  XM12
timestamp 1747747376
transform 1 0 7668 0 1 4228
box -278 -300 278 300
use sky130_fd_pr__nfet_g5v0d10v5_6XHUDR  XM13
timestamp 1747747376
transform 1 0 7668 0 1 4828
box -278 -300 278 300
use sky130_fd_pr__pfet_g5v0d10v5_6ELFTH  XM15
timestamp 1747747376
transform 1 0 5578 0 1 5695
box -308 -339 308 339
use sky130_fd_pr__nfet_g5v0d10v5_6XHUDR  XM16
timestamp 1747747376
transform 1 0 5256 0 1 4830
box -278 -300 278 300
use sky130_fd_pr__pfet_g5v0d10v5_6ELFTH  XM17
timestamp 1747747376
transform 1 0 4962 0 1 6373
box -308 -339 308 339
use sky130_fd_pr__pfet_g5v0d10v5_6ELFTH  XM18
timestamp 1747747376
transform 1 0 5578 0 1 6373
box -308 -339 308 339
use sky130_fd_pr__nfet_g5v0d10v5_6XHUDR  XM19
timestamp 1747747376
transform 1 0 5256 0 1 4230
box -278 -300 278 300
use sky130_fd_pr__nfet_g5v0d10v5_6XHUDR  XM20
timestamp 1747747376
transform 1 0 4700 0 1 4230
box -278 -300 278 300
use sky130_fd_pr__nfet_g5v0d10v5_6XHUDR  XM21
timestamp 1747747376
transform 1 0 1920 0 1 4230
box -278 -300 278 300
use sky130_fd_pr__pfet_g5v0d10v5_6ELFTH  XM22
timestamp 1747747376
transform 1 0 2498 0 1 6373
box -308 -339 308 339
use sky130_fd_pr__nfet_g5v0d10v5_6XHUDR  XM23
timestamp 1747747376
transform 1 0 1920 0 1 4828
box -278 -300 278 300
use sky130_fd_pr__pfet_g5v0d10v5_6ELFTH  XM24
timestamp 1747747376
transform 1 0 3114 0 1 6373
box -308 -339 308 339
use sky130_fd_pr__pfet_g5v0d10v5_6ELFTH  XM25
timestamp 1747747376
transform 1 0 3730 0 1 6373
box -308 -339 308 339
use sky130_fd_pr__pfet_g5v0d10v5_6ELFTH  XM26
timestamp 1747747376
transform 1 0 4346 0 1 6373
box -308 -339 308 339
use sky130_fd_pr__nfet_g5v0d10v5_6XHUDR  XM27
timestamp 1747747376
transform 1 0 4144 0 1 4230
box -278 -300 278 300
use sky130_fd_pr__nfet_g5v0d10v5_6XHUDR  XM28
timestamp 1747747376
transform 1 0 3588 0 1 4230
box -278 -300 278 300
use sky130_fd_pr__nfet_g5v0d10v5_6XHUDR  XM29
timestamp 1747747376
transform 1 0 3032 0 1 4230
box -278 -300 278 300
use sky130_fd_pr__nfet_g5v0d10v5_6XHUDR  XM30
timestamp 1747747376
transform 1 0 2476 0 1 4230
box -278 -300 278 300
use sky130_fd_pr__pfet_g5v0d10v5_6ELFTH  XM31
timestamp 1747747376
transform 1 0 6194 0 1 5695
box -308 -339 308 339
use sky130_fd_pr__nfet_g5v0d10v5_6XHUDR  XM32
timestamp 1747747376
transform 1 0 5812 0 1 4830
box -278 -300 278 300
use sky130_fd_pr__nfet_g5v0d10v5_6XHUDR  XM33
timestamp 1747747376
transform 1 0 1364 0 1 4828
box -278 -300 278 300
use sky130_fd_pr__pfet_g5v0d10v5_6ELFTH  XM34
timestamp 1747747376
transform 1 0 2498 0 1 5695
box -308 -339 308 339
use sky130_fd_pr__nfet_01v8_L7BSKG  XM35 paramcells
timestamp 1747747376
transform 1 0 10367 0 1 6113
box -211 -221 211 221
use sky130_fd_pr__nfet_g5v0d10v5_6XHUDR  XM36
timestamp 1747747376
transform 1 0 2476 0 1 4830
box -278 -300 278 300
use sky130_fd_pr__pfet_g5v0d10v5_6ELFTH  XM37
timestamp 1747747376
transform 1 0 6810 0 1 5695
box -308 -339 308 339
use sky130_fd_pr__nfet_g5v0d10v5_6XHUDR  XM38
timestamp 1747747376
transform 1 0 6368 0 1 4830
box -278 -300 278 300
use sky130_fd_pr__pfet_g5v0d10v5_6ELFTH  XM39
timestamp 1747747376
transform 1 0 6194 0 1 6373
box -308 -339 308 339
use sky130_fd_pr__pfet_g5v0d10v5_6ELFTH  XM40
timestamp 1747747376
transform 1 0 6810 0 1 6373
box -308 -339 308 339
use sky130_fd_pr__nfet_g5v0d10v5_6XHUDR  XM41
timestamp 1747747376
transform 1 0 6368 0 1 4230
box -278 -300 278 300
use sky130_fd_pr__nfet_g5v0d10v5_6XHUDR  XM42
timestamp 1747747376
transform 1 0 5812 0 1 4230
box -278 -300 278 300
<< labels >>
flabel metal2 12042 4786 12242 4986 0 FreeSans 256 0 0 0 ena
port 4 nsew
flabel metal2 12042 5630 12242 5830 0 FreeSans 256 0 0 0 dout
port 5 nsew
flabel metal1 12044 6364 12244 7121 0 FreeSans 256 0 0 0 dvss
port 2 nsew
flabel metal2 -24 7721 176 9715 0 FreeSans 256 0 0 0 avdd
port 0 nsew
flabel metal2 s 12144 7721 12244 9715 0 FreeSans 640 90 0 0 avdd
port 0 nsew
flabel metal1 12064 3634 12264 4391 0 FreeSans 256 0 0 0 dvdd
port 3 nsew
flabel metal2 -24 1050 176 3044 0 FreeSans 256 0 0 0 avss
port 1 nsew
flabel metal2 s 11934 1050 12242 3044 0 FreeSans 960 90 0 0 avss
port 1 nsew
<< properties >>
string FIXED_BBOX 0 0 12242 10724
<< end >>
